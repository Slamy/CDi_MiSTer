// verilator lint_off UNOPTFLAT
// verilator lint_off INITIALDLY
// verilator lint_off COMBDLY
// verilator lint_off CASEINCOMPLETE
// verilator lint_off UNSIGNED

module tg68k_alu_2_1_2_1
  (input  clk,
   input  reset,
   input  clkena_lw,
   input  [1:0] cpu,
   input  execopc,
   input  decodeopc,
   input  exe_condition,
   input  exec_tas,
   input  long_start,
   input  non_aligned,
   input  check_aligned,
   input  movem_presub,
   input  set_stop,
   input  z_error,
   input  [1:0] rot_bits,
   input  [88:0] exec,
   input  [31:0] op1out,
   input  [31:0] op2out,
   input  [31:0] reg_qa,
   input  [31:0] reg_qb,
   input  [15:0] opcode,
   input  [15:0] exe_opcode,
   input  [1:0] exe_datatype,
   input  [15:0] sndopc,
   input  [15:0] last_data_read,
   input  [15:0] data_read,
   input  [7:0] flagssr,
   input  [6:0] micro_state,
   input  [7:0] bf_ext_in,
   input  [5:0] bf_shift,
   input  [5:0] bf_width,
   input  [31:0] bf_ffo_offset,
   input  [4:0] bf_loffset,
   output [7:0] bf_ext_out,
   output set_v_flag,
   output [7:0] flags,
   output [2:0] c_out,
   output [31:0] addsub_q,
   output [31:0] aluout);
  wire [31:0] op1in;
  wire [31:0] addsub_a;
  wire [31:0] addsub_b;
  wire [33:0] notaddsub_b;
  wire [33:0] add_result;
  wire [2:0] addsub_ofl;
  wire opaddsub;
  wire [3:0] c_in;
  wire [2:0] flag_z;
  wire [3:0] set_flags;
  wire [7:0] ccrin;
  wire [3:0] last_flags1;
  wire [9:0] bcd_pur;
  wire [8:0] bcd_kor;
  wire halve_carry;
  wire vflag_a;
  wire bcd_a_carry;
  wire [8:0] bcd_a;
  wire [127:0] result_mulu;
  wire [63:0] result_div;
  wire [31:0] result_div_pre;
  wire set_mv_flag;
  wire v_flag;
  wire rot_rot;
  wire rot_x;
  wire rot_c;
  wire [31:0] rot_out;
  wire asl_vflag;
  wire [4:0] bit_number;
  wire [31:0] bits_out;
  wire one_bit_in;
  wire bchg;
  wire bset;
  wire [63:0] mulu_reg;
  wire [31:0] faktora;
  wire [31:0] faktorb;
  wire [63:0] div_reg;
  wire [63:0] div_quot;
  wire div_neg;
  wire div_bit;
  wire [32:0] div_sub;
  wire [32:0] div_over;
  wire nozero;
  wire div_qsign;
  wire [63:0] dividend;
  wire divs;
  wire signedop;
  wire op1_sign;
  wire [15:0] op2outext;
  wire [31:0] datareg;
  wire [31:0] bf_datareg;
  wire [39:0] result;
  wire [39:0] result_tmp;
  wire [31:0] unshifted_bitmask;
  wire [39:0] inmux0;
  wire [39:0] inmux1;
  wire [39:0] inmux2;
  wire [31:0] inmux3;
  wire [39:0] shifted_bitmask;
  wire [37:0] bitmaskmux0;
  wire [35:0] bitmaskmux1;
  wire [31:0] bitmaskmux2;
  wire [31:0] bitmaskmux3;
  wire [31:0] bf_set2;
  wire [39:0] shift;
  wire [5:0] bf_firstbit;
  wire [3:0] mux;
  wire [4:0] bitnr;
  wire [31:0] mask;
  wire mask_not_zero;
  wire bf_bset;
  wire bf_nflag;
  wire bf_bchg;
  wire bf_ins;
  wire bf_exts;
  wire bf_fffo;
  wire bf_d32;
  wire bf_s32;
  wire [33:0] hot_msb;
  wire [32:0] vector;
  wire [65:0] result_bs;
  wire [5:0] bit_nr;
  wire [5:0] bit_msb;
  wire [5:0] bs_shift;
  wire [5:0] bs_shift_mod;
  wire [32:0] asl_over;
  wire [32:0] asl_over_xor;
  wire [32:0] asr_sign;
  wire msb;
  wire [5:0] ring;
  wire [31:0] alu;
  wire [31:0] bsout;
  wire bs_v;
  wire bs_c;
  wire bs_x;
  wire n9938_o;
  wire n9939_o;
  wire [23:0] n9940_o;
  wire [6:0] n9941_o;
  wire n9942_o;
  wire [31:0] n9943_o;
  wire [31:0] n9944_o;
  wire [31:0] n9945_o;
  wire [31:0] n9946_o;
  wire [31:0] n9947_o;
  wire [31:0] n9948_o;
  wire n9949_o;
  wire n9950_o;
  wire n9951_o;
  wire [7:0] n9952_o;
  wire n9953_o;
  wire n9955_o;
  wire n9956_o;
  wire [31:0] n9957_o;
  wire [31:0] n9958_o;
  wire [31:0] n9959_o;
  wire n9960_o;
  wire n9962_o;
  wire n9963_o;
  wire n9965_o;
  wire [15:0] n9966_o;
  wire [15:0] n9967_o;
  wire [31:0] n9968_o;
  wire n9969_o;
  wire [31:0] n9970_o;
  wire [31:0] n9971_o;
  wire [31:0] n9972_o;
  wire [31:0] n9973_o;
  wire n9974_o;
  wire [31:0] n9975_o;
  wire n9976_o;
  wire [31:0] n9977_o;
  wire n9978_o;
  wire [3:0] n9979_o;
  wire [3:0] n9980_o;
  wire [7:0] n9981_o;
  wire n9982_o;
  wire [31:0] n9983_o;
  wire n9984_o;
  wire n9985_o;
  wire n9986_o;
  wire n9987_o;
  wire [15:0] n9988_o;
  wire [15:0] n9989_o;
  wire [31:0] n9990_o;
  wire n9991_o;
  wire n9992_o;
  wire n9993_o;
  wire n9994_o;
  wire [7:0] n9996_o;
  wire n9997_o;
  wire [3:0] n9998_o;
  wire [3:0] n9999_o;
  wire [7:0] n10000_o;
  wire [7:0] n10001_o;
  wire [7:0] n10002_o;
  wire [15:0] n10003_o;
  wire [7:0] n10004_o;
  wire [7:0] n10005_o;
  wire [7:0] n10006_o;
  wire [7:0] n10007_o;
  wire [7:0] n10008_o;
  wire [15:0] n10009_o;
  wire [15:0] n10010_o;
  wire [15:0] n10011_o;
  wire [15:0] n10012_o;
  wire [15:0] n10013_o;
  wire [15:0] n10014_o;
  wire [31:0] n10015_o;
  wire [31:0] n10016_o;
  wire [31:0] n10017_o;
  wire [31:0] n10018_o;
  wire [31:0] n10019_o;
  wire [31:0] n10020_o;
  wire [31:0] n10021_o;
  wire [7:0] n10022_o;
  wire [7:0] n10023_o;
  wire [23:0] n10024_o;
  wire [23:0] n10025_o;
  wire [23:0] n10026_o;
  wire [31:0] n10027_o;
  wire [31:0] n10028_o;
  wire [31:0] n10029_o;
  wire [31:0] n10030_o;
  wire [31:0] n10031_o;
  wire [7:0] n10032_o;
  wire [7:0] n10033_o;
  wire [23:0] n10034_o;
  wire [23:0] n10035_o;
  wire [23:0] n10036_o;
  wire n10041_o;
  wire n10042_o;
  wire n10043_o;
  wire n10044_o;
  wire [1:0] n10045_o;
  wire n10046_o;
  wire [2:0] n10047_o;
  wire [28:0] n10048_o;
  wire [31:0] n10049_o;
  wire [1:0] n10050_o;
  wire [31:0] n10052_o;
  wire [31:0] n10053_o;
  wire [31:0] n10054_o;
  wire n10055_o;
  wire n10058_o;
  wire n10060_o;
  wire [3:0] n10061_o;
  wire [7:0] n10063_o;
  wire [11:0] n10065_o;
  wire [3:0] n10066_o;
  wire [15:0] n10067_o;
  wire n10068_o;
  wire n10069_o;
  wire n10070_o;
  wire n10071_o;
  wire n10072_o;
  wire n10073_o;
  wire n10074_o;
  wire n10075_o;
  wire n10077_o;
  wire n10078_o;
  wire n10079_o;
  wire n10080_o;
  wire n10081_o;
  wire n10082_o;
  wire n10084_o;
  wire n10085_o;
  wire n10086_o;
  wire n10087_o;
  wire n10088_o;
  wire n10089_o;
  wire n10090_o;
  wire n10091_o;
  wire [31:0] n10094_o;
  wire [31:0] n10096_o;
  wire [31:0] n10098_o;
  wire n10099_o;
  wire n10100_o;
  wire n10101_o;
  wire n10102_o;
  wire n10103_o;
  wire n10105_o;
  wire n10106_o;
  wire [31:0] n10107_o;
  wire n10108_o;
  wire n10109_o;
  wire [15:0] n10110_o;
  wire [15:0] n10111_o;
  wire [15:0] n10112_o;
  wire [15:0] n10113_o;
  wire [15:0] n10114_o;
  wire n10116_o;
  wire n10117_o;
  wire n10118_o;
  wire n10119_o;
  wire n10120_o;
  wire n10121_o;
  wire n10122_o;
  wire [31:0] n10124_o;
  wire [31:0] n10125_o;
  wire n10126_o;
  wire n10127_o;
  wire n10129_o;
  wire [31:0] n10132_o;
  wire [31:0] n10133_o;
  wire [31:0] n10134_o;
  wire [31:0] n10135_o;
  wire [31:0] n10136_o;
  wire [31:0] n10137_o;
  wire n10138_o;
  wire n10139_o;
  wire [32:0] n10141_o;
  wire n10142_o;
  wire [33:0] n10143_o;
  wire [32:0] n10145_o;
  wire n10146_o;
  wire [33:0] n10147_o;
  wire [33:0] n10148_o;
  wire [33:0] n10149_o;
  wire [32:0] n10151_o;
  wire n10152_o;
  wire [33:0] n10153_o;
  wire [33:0] n10154_o;
  wire n10155_o;
  wire n10156_o;
  wire n10157_o;
  wire n10158_o;
  wire n10159_o;
  wire n10160_o;
  wire n10161_o;
  wire n10162_o;
  wire n10163_o;
  wire n10164_o;
  wire n10165_o;
  wire [31:0] n10166_o;
  wire n10167_o;
  wire n10168_o;
  wire n10169_o;
  wire n10170_o;
  wire n10171_o;
  wire n10172_o;
  wire n10173_o;
  wire n10174_o;
  wire n10175_o;
  wire n10176_o;
  wire n10177_o;
  wire n10178_o;
  wire n10179_o;
  wire n10180_o;
  wire n10181_o;
  wire n10182_o;
  wire n10183_o;
  wire n10184_o;
  wire n10185_o;
  wire n10186_o;
  wire n10187_o;
  wire [2:0] n10188_o;
  wire n10192_o;
  wire [8:0] n10193_o;
  wire [9:0] n10194_o;
  wire n10195_o;
  wire n10196_o;
  wire n10197_o;
  wire n10198_o;
  wire n10199_o;
  wire [3:0] n10202_o;
  localparam [8:0] n10203_o = 9'b000000000;
  wire n10205_o;
  wire [3:0] n10207_o;
  wire [3:0] n10208_o;
  wire n10209_o;
  wire n10210_o;
  wire n10211_o;
  wire n10212_o;
  wire n10213_o;
  wire n10214_o;
  wire [8:0] n10215_o;
  wire [8:0] n10216_o;
  wire n10217_o;
  wire n10218_o;
  wire n10219_o;
  wire n10220_o;
  wire n10221_o;
  wire [3:0] n10223_o;
  wire n10224_o;
  wire n10225_o;
  wire n10226_o;
  wire n10227_o;
  wire n10228_o;
  wire n10229_o;
  wire n10230_o;
  wire n10231_o;
  wire n10232_o;
  wire n10233_o;
  wire n10234_o;
  wire n10235_o;
  wire n10236_o;
  wire [3:0] n10238_o;
  wire n10239_o;
  wire n10240_o;
  wire n10241_o;
  wire n10242_o;
  wire [8:0] n10243_o;
  wire [8:0] n10244_o;
  wire [7:0] n10245_o;
  wire [7:0] n10246_o;
  wire [7:0] n10247_o;
  wire n10248_o;
  wire [8:0] n10249_o;
  wire n10250_o;
  wire n10252_o;
  wire n10253_o;
  wire n10254_o;
  wire n10255_o;
  wire [1:0] n10260_o;
  wire n10262_o;
  wire n10264_o;
  wire [1:0] n10265_o;
  reg n10268_o;
  reg n10272_o;
  wire n10278_o;
  wire n10279_o;
  wire [1:0] n10280_o;
  wire n10282_o;
  wire [4:0] n10283_o;
  wire [2:0] n10284_o;
  wire [4:0] n10286_o;
  wire [4:0] n10287_o;
  wire [1:0] n10288_o;
  wire n10290_o;
  wire [4:0] n10291_o;
  wire [2:0] n10292_o;
  wire [4:0] n10294_o;
  wire [4:0] n10295_o;
  wire [4:0] n10296_o;
  wire n10302_o;
  wire n10303_o;
  wire n10304_o;
  wire [1:0] n10310_o;
  wire n10312_o;
  wire n10315_o;
  wire [2:0] n10317_o;
  wire n10319_o;
  wire n10321_o;
  wire n10323_o;
  wire n10325_o;
  wire n10327_o;
  wire [4:0] n10328_o;
  reg n10331_o;
  reg n10335_o;
  reg n10339_o;
  reg n10343_o;
  reg n10347_o;
  reg n10350_o;
  wire [1:0] n10351_o;
  wire n10353_o;
  wire n10356_o;
  wire [7:0] n10358_o;
  wire [4:0] n10376_o;
  wire n10378_o;
  wire n10381_o;
  wire n10382_o;
  wire n10383_o;
  wire n10384_o;
  wire n10389_o;
  localparam [31:0] n10390_o = 32'b00000000000000000000000000000000;
  wire [4:0] n10392_o;
  wire n10394_o;
  wire n10397_o;
  wire n10398_o;
  wire n10399_o;
  wire n10400_o;
  wire n10404_o;
  wire n10405_o;
  wire [4:0] n10407_o;
  wire n10409_o;
  wire n10412_o;
  wire n10413_o;
  wire n10414_o;
  wire n10415_o;
  wire n10419_o;
  wire n10420_o;
  wire [4:0] n10422_o;
  wire n10424_o;
  wire n10427_o;
  wire n10428_o;
  wire n10429_o;
  wire n10430_o;
  wire n10434_o;
  wire n10435_o;
  wire [4:0] n10437_o;
  wire n10439_o;
  wire n10442_o;
  wire n10443_o;
  wire n10444_o;
  wire n10445_o;
  wire n10449_o;
  wire n10450_o;
  wire [4:0] n10452_o;
  wire n10454_o;
  wire n10457_o;
  wire n10458_o;
  wire n10459_o;
  wire n10460_o;
  wire n10464_o;
  wire n10465_o;
  wire [4:0] n10467_o;
  wire n10469_o;
  wire n10472_o;
  wire n10473_o;
  wire n10474_o;
  wire n10475_o;
  wire n10479_o;
  wire n10480_o;
  wire [4:0] n10482_o;
  wire n10484_o;
  wire n10487_o;
  wire n10488_o;
  wire n10489_o;
  wire n10490_o;
  wire n10494_o;
  wire n10495_o;
  wire [4:0] n10497_o;
  wire n10499_o;
  wire n10502_o;
  wire n10503_o;
  wire n10504_o;
  wire n10505_o;
  wire n10509_o;
  wire n10510_o;
  wire [4:0] n10512_o;
  wire n10514_o;
  wire n10517_o;
  wire n10518_o;
  wire n10519_o;
  wire n10520_o;
  wire n10524_o;
  wire n10525_o;
  wire [4:0] n10527_o;
  wire n10529_o;
  wire n10532_o;
  wire n10533_o;
  wire n10534_o;
  wire n10535_o;
  wire n10539_o;
  wire n10540_o;
  wire [4:0] n10542_o;
  wire n10544_o;
  wire n10547_o;
  wire n10548_o;
  wire n10549_o;
  wire n10550_o;
  wire n10554_o;
  wire n10555_o;
  wire [4:0] n10557_o;
  wire n10559_o;
  wire n10562_o;
  wire n10563_o;
  wire n10564_o;
  wire n10565_o;
  wire n10569_o;
  wire n10570_o;
  wire [4:0] n10572_o;
  wire n10574_o;
  wire n10577_o;
  wire n10578_o;
  wire n10579_o;
  wire n10580_o;
  wire n10584_o;
  wire n10585_o;
  wire [4:0] n10587_o;
  wire n10589_o;
  wire n10592_o;
  wire n10593_o;
  wire n10594_o;
  wire n10595_o;
  wire n10599_o;
  wire n10600_o;
  wire [4:0] n10602_o;
  wire n10604_o;
  wire n10607_o;
  wire n10608_o;
  wire n10609_o;
  wire n10610_o;
  wire n10614_o;
  wire n10615_o;
  wire [4:0] n10617_o;
  wire n10619_o;
  wire n10622_o;
  wire n10623_o;
  wire n10624_o;
  wire n10625_o;
  wire n10629_o;
  wire n10630_o;
  wire [4:0] n10632_o;
  wire n10634_o;
  wire n10637_o;
  wire n10638_o;
  wire n10639_o;
  wire n10640_o;
  wire n10644_o;
  wire n10645_o;
  wire [4:0] n10647_o;
  wire n10649_o;
  wire n10652_o;
  wire n10653_o;
  wire n10654_o;
  wire n10655_o;
  wire n10659_o;
  wire n10660_o;
  wire [4:0] n10662_o;
  wire n10664_o;
  wire n10667_o;
  wire n10668_o;
  wire n10669_o;
  wire n10670_o;
  wire n10674_o;
  wire n10675_o;
  wire [4:0] n10677_o;
  wire n10679_o;
  wire n10682_o;
  wire n10683_o;
  wire n10684_o;
  wire n10685_o;
  wire n10689_o;
  wire n10690_o;
  wire [4:0] n10692_o;
  wire n10694_o;
  wire n10697_o;
  wire n10698_o;
  wire n10699_o;
  wire n10700_o;
  wire n10704_o;
  wire n10705_o;
  wire [4:0] n10707_o;
  wire n10709_o;
  wire n10712_o;
  wire n10713_o;
  wire n10714_o;
  wire n10715_o;
  wire n10719_o;
  wire n10720_o;
  wire [4:0] n10722_o;
  wire n10724_o;
  wire n10727_o;
  wire n10728_o;
  wire n10729_o;
  wire n10730_o;
  wire n10734_o;
  wire n10735_o;
  wire [4:0] n10737_o;
  wire n10739_o;
  wire n10742_o;
  wire n10743_o;
  wire n10744_o;
  wire n10745_o;
  wire n10749_o;
  wire n10750_o;
  wire [4:0] n10752_o;
  wire n10754_o;
  wire n10757_o;
  wire n10758_o;
  wire n10759_o;
  wire n10760_o;
  wire n10764_o;
  wire n10765_o;
  wire [4:0] n10767_o;
  wire n10769_o;
  wire n10772_o;
  wire n10773_o;
  wire n10774_o;
  wire n10775_o;
  wire n10779_o;
  wire n10780_o;
  wire [4:0] n10782_o;
  wire n10784_o;
  wire n10787_o;
  wire n10788_o;
  wire n10789_o;
  wire n10790_o;
  wire n10794_o;
  wire n10795_o;
  wire [4:0] n10797_o;
  wire n10799_o;
  wire n10802_o;
  wire n10803_o;
  wire n10804_o;
  wire n10805_o;
  wire n10809_o;
  wire n10810_o;
  wire [4:0] n10812_o;
  wire n10814_o;
  wire n10817_o;
  wire n10818_o;
  wire n10819_o;
  wire n10820_o;
  wire n10824_o;
  wire n10825_o;
  wire [4:0] n10827_o;
  wire n10829_o;
  wire n10832_o;
  wire n10833_o;
  wire n10834_o;
  wire n10835_o;
  wire n10836_o;
  wire n10837_o;
  wire n10838_o;
  wire n10839_o;
  wire n10840_o;
  wire n10841_o;
  wire [4:0] n10842_o;
  wire n10844_o;
  wire n10847_o;
  wire n10848_o;
  wire [4:0] n10850_o;
  wire n10853_o;
  wire [31:0] n10854_o;
  wire [31:0] n10855_o;
  wire n10856_o;
  wire [15:0] n10857_o;
  wire [15:0] n10858_o;
  wire [31:0] n10859_o;
  wire [31:0] n10860_o;
  wire n10861_o;
  wire [23:0] n10862_o;
  wire [7:0] n10863_o;
  wire [31:0] n10864_o;
  wire [31:0] n10865_o;
  wire n10866_o;
  wire [35:0] n10868_o;
  wire [3:0] n10869_o;
  wire [3:0] n10870_o;
  wire [3:0] n10871_o;
  wire [31:0] n10872_o;
  wire [35:0] n10874_o;
  wire [35:0] n10875_o;
  wire [35:0] n10876_o;
  wire n10877_o;
  wire [37:0] n10879_o;
  wire [1:0] n10880_o;
  wire [1:0] n10881_o;
  wire [1:0] n10882_o;
  wire [35:0] n10883_o;
  wire [37:0] n10885_o;
  wire [37:0] n10886_o;
  wire [37:0] n10887_o;
  wire n10888_o;
  wire [38:0] n10890_o;
  wire [39:0] n10892_o;
  wire n10893_o;
  wire n10894_o;
  wire n10895_o;
  wire [38:0] n10896_o;
  wire [39:0] n10898_o;
  wire [39:0] n10899_o;
  wire [39:0] n10900_o;
  wire [39:0] n10901_o;
  wire [7:0] n10902_o;
  wire [7:0] n10903_o;
  wire [7:0] n10904_o;
  wire [31:0] n10905_o;
  wire n10906_o;
  wire n10907_o;
  wire [38:0] n10908_o;
  wire [39:0] n10909_o;
  wire [39:0] n10910_o;
  wire n10911_o;
  wire [1:0] n10912_o;
  wire [37:0] n10913_o;
  wire [39:0] n10914_o;
  wire [39:0] n10915_o;
  wire n10916_o;
  wire [3:0] n10917_o;
  wire [35:0] n10918_o;
  wire [39:0] n10919_o;
  wire [39:0] n10920_o;
  wire n10921_o;
  wire [7:0] n10922_o;
  wire [23:0] n10923_o;
  wire [31:0] n10924_o;
  wire [31:0] n10925_o;
  wire [31:0] n10926_o;
  wire n10927_o;
  wire [15:0] n10928_o;
  wire [15:0] n10929_o;
  wire [31:0] n10930_o;
  wire [31:0] n10931_o;
  wire [7:0] n10932_o;
  wire [31:0] n10933_o;
  wire [7:0] n10934_o;
  wire [39:0] n10935_o;
  localparam [39:0] n10936_o = 40'b0000000000000000000000000000000000000000;
  wire [39:0] n10938_o;
  localparam [39:0] n10940_o = 40'b1111111111111111111111111111111111111111;
  wire [39:0] n10942_o;
  wire [39:0] n10943_o;
  wire [39:0] n10944_o;
  wire n10945_o;
  wire n10946_o;
  wire n10947_o;
  wire n10948_o;
  wire n10949_o;
  wire n10950_o;
  wire n10951_o;
  wire n10952_o;
  wire n10953_o;
  wire n10954_o;
  wire n10962_o;
  wire n10963_o;
  wire n10964_o;
  wire n10965_o;
  wire n10966_o;
  wire n10967_o;
  wire n10968_o;
  wire n10969_o;
  wire n10970_o;
  wire n10971_o;
  wire n10979_o;
  wire n10980_o;
  wire n10981_o;
  wire n10982_o;
  wire n10983_o;
  wire n10984_o;
  wire n10985_o;
  wire n10986_o;
  wire n10987_o;
  wire n10988_o;
  wire n10996_o;
  wire n10997_o;
  wire n10998_o;
  wire n10999_o;
  wire n11000_o;
  wire n11001_o;
  wire n11002_o;
  wire n11003_o;
  wire n11004_o;
  wire n11005_o;
  wire n11013_o;
  wire n11014_o;
  wire n11015_o;
  wire n11016_o;
  wire n11017_o;
  wire n11018_o;
  wire n11019_o;
  wire n11020_o;
  wire n11021_o;
  wire n11022_o;
  wire n11030_o;
  wire n11031_o;
  wire n11032_o;
  wire n11033_o;
  wire n11034_o;
  wire n11035_o;
  wire n11036_o;
  wire n11037_o;
  wire n11038_o;
  wire n11039_o;
  wire n11047_o;
  wire n11048_o;
  wire n11049_o;
  wire n11050_o;
  wire n11051_o;
  wire n11052_o;
  wire n11053_o;
  wire n11054_o;
  wire n11055_o;
  wire n11056_o;
  wire n11064_o;
  wire n11065_o;
  wire n11066_o;
  wire n11067_o;
  wire n11068_o;
  wire n11069_o;
  wire n11070_o;
  wire n11071_o;
  wire n11072_o;
  wire n11073_o;
  wire n11081_o;
  wire n11082_o;
  wire n11083_o;
  wire n11084_o;
  wire n11085_o;
  wire n11086_o;
  wire n11087_o;
  wire n11088_o;
  wire n11089_o;
  wire n11090_o;
  wire n11098_o;
  wire n11099_o;
  wire n11100_o;
  wire n11101_o;
  wire n11102_o;
  wire n11103_o;
  wire n11104_o;
  wire n11105_o;
  wire n11106_o;
  wire n11107_o;
  wire n11115_o;
  wire n11116_o;
  wire n11117_o;
  wire n11118_o;
  wire n11119_o;
  wire n11120_o;
  wire n11121_o;
  wire n11122_o;
  wire n11123_o;
  wire n11124_o;
  wire n11132_o;
  wire n11133_o;
  wire n11134_o;
  wire n11135_o;
  wire n11136_o;
  wire n11137_o;
  wire n11138_o;
  wire n11139_o;
  wire n11140_o;
  wire n11141_o;
  wire n11149_o;
  wire n11150_o;
  wire n11151_o;
  wire n11152_o;
  wire n11153_o;
  wire n11154_o;
  wire n11155_o;
  wire n11156_o;
  wire n11157_o;
  wire n11158_o;
  wire n11166_o;
  wire n11167_o;
  wire n11168_o;
  wire n11169_o;
  wire n11170_o;
  wire n11171_o;
  wire n11172_o;
  wire n11173_o;
  wire n11174_o;
  wire n11175_o;
  wire n11183_o;
  wire n11184_o;
  wire n11185_o;
  wire n11186_o;
  wire n11187_o;
  wire n11188_o;
  wire n11189_o;
  wire n11190_o;
  wire n11191_o;
  wire n11192_o;
  wire n11200_o;
  wire n11201_o;
  wire n11202_o;
  wire n11203_o;
  wire n11204_o;
  wire n11205_o;
  wire n11206_o;
  wire n11207_o;
  wire n11208_o;
  wire n11209_o;
  wire n11217_o;
  wire n11218_o;
  wire n11219_o;
  wire n11220_o;
  wire n11221_o;
  wire n11222_o;
  wire n11223_o;
  wire n11224_o;
  wire n11225_o;
  wire n11226_o;
  wire n11234_o;
  wire n11235_o;
  wire n11236_o;
  wire n11237_o;
  wire n11238_o;
  wire n11239_o;
  wire n11240_o;
  wire n11241_o;
  wire n11242_o;
  wire n11243_o;
  wire n11251_o;
  wire n11252_o;
  wire n11253_o;
  wire n11254_o;
  wire n11255_o;
  wire n11256_o;
  wire n11257_o;
  wire n11258_o;
  wire n11259_o;
  wire n11260_o;
  wire n11268_o;
  wire n11269_o;
  wire n11270_o;
  wire n11271_o;
  wire n11272_o;
  wire n11273_o;
  wire n11274_o;
  wire n11275_o;
  wire n11276_o;
  wire n11277_o;
  wire n11285_o;
  wire n11286_o;
  wire n11287_o;
  wire n11288_o;
  wire n11289_o;
  wire n11290_o;
  wire n11291_o;
  wire n11292_o;
  wire n11293_o;
  wire n11294_o;
  wire n11302_o;
  wire n11303_o;
  wire n11304_o;
  wire n11305_o;
  wire n11306_o;
  wire n11307_o;
  wire n11308_o;
  wire n11309_o;
  wire n11310_o;
  wire n11311_o;
  wire n11319_o;
  wire n11320_o;
  wire n11321_o;
  wire n11322_o;
  wire n11323_o;
  wire n11324_o;
  wire n11325_o;
  wire n11326_o;
  wire n11327_o;
  wire n11328_o;
  wire n11336_o;
  wire n11337_o;
  wire n11338_o;
  wire n11339_o;
  wire n11340_o;
  wire n11341_o;
  wire n11342_o;
  wire n11343_o;
  wire n11344_o;
  wire n11345_o;
  wire n11353_o;
  wire n11354_o;
  wire n11355_o;
  wire n11356_o;
  wire n11357_o;
  wire n11358_o;
  wire n11359_o;
  wire n11360_o;
  wire n11361_o;
  wire n11362_o;
  wire n11370_o;
  wire n11371_o;
  wire n11372_o;
  wire n11373_o;
  wire n11374_o;
  wire n11375_o;
  wire n11376_o;
  wire n11377_o;
  wire n11378_o;
  wire n11379_o;
  wire n11387_o;
  wire n11388_o;
  wire n11389_o;
  wire n11390_o;
  wire n11391_o;
  wire n11392_o;
  wire n11393_o;
  wire n11394_o;
  wire n11395_o;
  wire n11396_o;
  wire n11404_o;
  wire n11405_o;
  wire n11406_o;
  wire n11407_o;
  wire n11408_o;
  wire n11409_o;
  wire n11410_o;
  wire n11411_o;
  wire n11412_o;
  wire n11413_o;
  wire n11421_o;
  wire n11422_o;
  wire n11423_o;
  wire n11424_o;
  wire n11425_o;
  wire n11426_o;
  wire n11427_o;
  wire n11428_o;
  wire n11429_o;
  wire n11430_o;
  wire n11438_o;
  wire n11439_o;
  wire n11440_o;
  wire n11441_o;
  wire n11442_o;
  wire n11443_o;
  wire n11444_o;
  wire n11445_o;
  wire n11446_o;
  wire n11447_o;
  wire n11455_o;
  wire n11456_o;
  wire n11457_o;
  wire n11458_o;
  wire n11459_o;
  wire n11460_o;
  wire n11461_o;
  wire n11462_o;
  wire n11463_o;
  wire n11464_o;
  wire n11472_o;
  wire n11473_o;
  wire n11474_o;
  wire n11475_o;
  wire n11476_o;
  wire n11477_o;
  wire n11478_o;
  wire n11479_o;
  wire n11480_o;
  wire n11481_o;
  wire n11489_o;
  wire n11490_o;
  wire n11491_o;
  wire n11492_o;
  wire n11493_o;
  wire n11494_o;
  wire n11495_o;
  wire n11496_o;
  wire n11497_o;
  wire n11498_o;
  wire n11506_o;
  wire n11507_o;
  wire n11508_o;
  wire n11509_o;
  wire n11510_o;
  wire n11511_o;
  wire n11512_o;
  wire n11513_o;
  wire n11514_o;
  wire n11515_o;
  wire n11523_o;
  wire n11524_o;
  wire n11525_o;
  wire n11526_o;
  wire n11527_o;
  wire n11528_o;
  wire n11529_o;
  wire n11530_o;
  wire n11531_o;
  wire n11532_o;
  wire n11540_o;
  wire n11541_o;
  wire n11542_o;
  wire n11543_o;
  wire n11544_o;
  wire n11545_o;
  wire n11546_o;
  wire n11547_o;
  wire n11548_o;
  wire n11549_o;
  wire n11557_o;
  wire n11558_o;
  wire n11559_o;
  wire n11560_o;
  wire n11561_o;
  wire n11562_o;
  wire n11563_o;
  wire n11564_o;
  wire n11565_o;
  wire n11566_o;
  wire n11574_o;
  wire n11575_o;
  wire n11576_o;
  wire n11577_o;
  wire n11578_o;
  wire n11579_o;
  wire n11580_o;
  wire n11581_o;
  wire n11582_o;
  wire n11583_o;
  wire n11591_o;
  wire n11592_o;
  wire n11593_o;
  wire n11594_o;
  wire n11595_o;
  wire n11596_o;
  wire n11597_o;
  wire n11598_o;
  wire n11599_o;
  wire n11600_o;
  wire n11601_o;
  wire n11602_o;
  wire n11603_o;
  wire n11604_o;
  wire n11605_o;
  wire n11606_o;
  wire n11607_o;
  wire n11608_o;
  wire n11609_o;
  wire n11610_o;
  wire [5:0] n11612_o;
  wire [5:0] n11613_o;
  wire [5:0] n11614_o;
  wire [3:0] n11615_o;
  wire n11617_o;
  wire [3:0] n11618_o;
  wire n11620_o;
  wire [3:0] n11621_o;
  wire n11623_o;
  wire [3:0] n11624_o;
  wire n11626_o;
  wire [3:0] n11628_o;
  wire n11630_o;
  wire [3:0] n11631_o;
  wire n11633_o;
  wire [3:0] n11635_o;
  wire n11637_o;
  wire [3:0] n11639_o;
  wire [3:0] n11640_o;
  wire [3:0] n11641_o;
  wire n11643_o;
  wire [3:0] n11644_o;
  wire [3:0] n11646_o;
  wire [1:0] n11647_o;
  wire n11648_o;
  wire n11649_o;
  wire n11650_o;
  wire n11652_o;
  wire [3:0] n11653_o;
  wire [3:0] n11654_o;
  wire [1:0] n11655_o;
  wire [1:0] n11657_o;
  wire [3:0] n11658_o;
  wire [3:0] n11661_o;
  wire [1:0] n11662_o;
  wire [2:0] n11663_o;
  wire [1:0] n11664_o;
  wire [1:0] n11665_o;
  wire n11666_o;
  wire n11668_o;
  wire [3:0] n11669_o;
  wire [3:0] n11671_o;
  wire [2:0] n11672_o;
  wire n11673_o;
  wire n11675_o;
  wire n11676_o;
  wire n11677_o;
  wire n11678_o;
  wire n11680_o;
  wire [3:0] n11681_o;
  wire [3:0] n11683_o;
  wire [2:0] n11684_o;
  wire n11685_o;
  wire n11686_o;
  wire [1:0] n11687_o;
  wire [1:0] n11689_o;
  wire [3:0] n11690_o;
  wire [3:0] n11691_o;
  wire [2:0] n11692_o;
  wire [2:0] n11694_o;
  localparam [4:0] n11695_o = 5'b11111;
  wire [1:0] n11697_o;
  wire n11699_o;
  wire n11701_o;
  wire n11702_o;
  wire n11704_o;
  wire n11705_o;
  wire n11708_o;
  wire n11709_o;
  wire n11710_o;
  wire n11712_o;
  wire n11713_o;
  wire n11714_o;
  wire n11716_o;
  wire n11717_o;
  wire [1:0] n11718_o;
  wire n11719_o;
  wire n11720_o;
  wire n11721_o;
  wire n11722_o;
  wire n11723_o;
  wire n11726_o;
  wire [1:0] n11731_o;
  wire n11732_o;
  wire n11734_o;
  wire n11735_o;
  wire n11737_o;
  wire n11739_o;
  wire n11740_o;
  wire n11741_o;
  wire n11743_o;
  wire [2:0] n11744_o;
  reg n11745_o;
  wire n11763_o;
  wire n11764_o;
  wire n11766_o;
  wire n11767_o;
  wire n11769_o;
  wire n11770_o;
  wire n11773_o;
  wire n11774_o;
  wire n11794_o;
  wire n11795_o;
  wire n11798_o;
  wire n11799_o;
  wire [31:0] n11800_o;
  wire n11805_o;
  wire [1:0] n11806_o;
  wire n11808_o;
  wire n11810_o;
  wire n11812_o;
  wire n11813_o;
  wire n11815_o;
  wire [2:0] n11816_o;
  reg [5:0] n11821_o;
  wire [1:0] n11822_o;
  wire n11824_o;
  wire n11826_o;
  wire n11828_o;
  wire n11829_o;
  wire n11831_o;
  wire [2:0] n11832_o;
  reg [5:0] n11837_o;
  wire [5:0] n11838_o;
  wire [1:0] n11840_o;
  wire n11842_o;
  wire n11843_o;
  wire n11844_o;
  wire n11845_o;
  wire n11846_o;
  wire [5:0] n11847_o;
  wire [2:0] n11848_o;
  wire [2:0] n11849_o;
  wire n11851_o;
  wire [2:0] n11854_o;
  wire [5:0] n11855_o;
  wire [5:0] n11856_o;
  wire [5:0] n11858_o;
  localparam [33:0] n11861_o = 34'b0000000000000000000000000000000000;
  wire n11865_o;
  wire [5:0] n11866_o;
  wire [5:0] n11868_o;
  wire [30:0] n11870_o;
  wire [31:0] n11872_o;
  wire [30:0] n11873_o;
  wire [31:0] n11875_o;
  wire [31:0] n11876_o;
  wire [32:0] n11877_o;
  wire [1:0] n11878_o;
  wire n11881_o;
  wire n11884_o;
  wire n11886_o;
  wire n11887_o;
  wire [1:0] n11888_o;
  wire n11889_o;
  reg n11890_o;
  wire n11891_o;
  reg n11892_o;
  wire [7:0] n11894_o;
  wire [15:0] n11895_o;
  wire [6:0] n11896_o;
  wire [31:0] n11897_o;
  wire [32:0] n11899_o;
  wire [32:0] n11900_o;
  wire n11902_o;
  wire n11903_o;
  wire n11904_o;
  wire n11905_o;
  wire n11906_o;
  wire n11908_o;
  wire n11910_o;
  wire n11911_o;
  wire n11912_o;
  wire [1:0] n11913_o;
  wire n11914_o;
  wire n11916_o;
  wire n11917_o;
  wire n11919_o;
  wire n11921_o;
  wire n11922_o;
  wire n11923_o;
  wire n11925_o;
  wire [2:0] n11926_o;
  reg n11927_o;
  wire n11928_o;
  wire n11930_o;
  wire n11931_o;
  wire [1:0] n11932_o;
  wire [7:0] n11933_o;
  wire [7:0] n11934_o;
  wire [7:0] n11935_o;
  wire n11936_o;
  wire n11938_o;
  wire [15:0] n11939_o;
  wire [15:0] n11940_o;
  wire [15:0] n11941_o;
  wire n11942_o;
  wire n11944_o;
  wire n11946_o;
  wire n11947_o;
  wire [31:0] n11948_o;
  wire [31:0] n11949_o;
  wire [31:0] n11950_o;
  wire n11951_o;
  wire n11953_o;
  wire [2:0] n11954_o;
  wire [7:0] n11955_o;
  wire [7:0] n11956_o;
  reg [7:0] n11958_o;
  wire [7:0] n11959_o;
  wire [7:0] n11960_o;
  reg [7:0] n11962_o;
  wire [15:0] n11963_o;
  reg [15:0] n11965_o;
  reg n11966_o;
  wire n11967_o;
  wire n11968_o;
  wire n11969_o;
  wire n11971_o;
  wire [1:0] n11972_o;
  wire [7:0] n11973_o;
  wire [7:0] n11974_o;
  wire [7:0] n11975_o;
  wire n11976_o;
  wire n11977_o;
  wire n11978_o;
  wire n11980_o;
  wire [15:0] n11981_o;
  wire [15:0] n11982_o;
  wire [15:0] n11983_o;
  wire n11984_o;
  wire n11985_o;
  wire n11986_o;
  wire n11988_o;
  wire n11990_o;
  wire n11991_o;
  wire [31:0] n11992_o;
  wire [31:0] n11993_o;
  wire [31:0] n11994_o;
  wire n11995_o;
  wire n11996_o;
  wire n11997_o;
  wire n11999_o;
  wire [2:0] n12000_o;
  wire [7:0] n12001_o;
  wire [7:0] n12002_o;
  reg [7:0] n12004_o;
  wire [7:0] n12005_o;
  wire [7:0] n12006_o;
  reg [7:0] n12008_o;
  wire [15:0] n12009_o;
  reg [15:0] n12011_o;
  reg n12012_o;
  wire n12013_o;
  wire n12014_o;
  wire [31:0] n12015_o;
  wire [31:0] n12016_o;
  wire [31:0] n12017_o;
  wire [31:0] n12018_o;
  wire [31:0] n12019_o;
  wire n12020_o;
  wire [31:0] n12021_o;
  wire [31:0] n12022_o;
  wire n12024_o;
  wire n12025_o;
  wire n12027_o;
  wire n12029_o;
  wire n12030_o;
  wire n12032_o;
  wire n12033_o;
  wire n12035_o;
  wire n12036_o;
  wire n12037_o;
  wire n12039_o;
  wire n12041_o;
  wire [5:0] n12043_o;
  wire n12045_o;
  wire [5:0] n12047_o;
  wire n12049_o;
  wire [5:0] n12051_o;
  wire n12053_o;
  wire [5:0] n12055_o;
  wire n12057_o;
  wire [5:0] n12059_o;
  wire n12061_o;
  wire [5:0] n12063_o;
  wire [5:0] n12064_o;
  wire [5:0] n12065_o;
  wire [5:0] n12066_o;
  wire [5:0] n12067_o;
  wire [5:0] n12068_o;
  wire [5:0] n12069_o;
  wire [5:0] n12071_o;
  wire n12073_o;
  wire n12075_o;
  wire [5:0] n12077_o;
  wire n12079_o;
  wire [5:0] n12081_o;
  wire n12083_o;
  wire [5:0] n12085_o;
  wire [5:0] n12086_o;
  wire [5:0] n12087_o;
  wire [5:0] n12088_o;
  wire n12090_o;
  wire n12092_o;
  wire [5:0] n12094_o;
  wire [5:0] n12095_o;
  wire n12097_o;
  wire [2:0] n12098_o;
  wire [5:0] n12100_o;
  wire n12102_o;
  wire [3:0] n12103_o;
  wire [5:0] n12105_o;
  wire n12107_o;
  wire [4:0] n12108_o;
  wire [5:0] n12110_o;
  wire n12112_o;
  wire [5:0] n12113_o;
  reg [5:0] n12115_o;
  wire n12116_o;
  wire n12117_o;
  wire [5:0] n12118_o;
  wire [5:0] n12119_o;
  wire n12120_o;
  wire n12121_o;
  wire n12122_o;
  wire n12123_o;
  wire [5:0] n12125_o;
  wire [5:0] n12126_o;
  wire n12127_o;
  wire n12128_o;
  wire n12129_o;
  wire [5:0] n12131_o;
  wire [5:0] n12132_o;
  wire [5:0] n12133_o;
  wire n12134_o;
  wire n12135_o;
  wire n12136_o;
  wire [5:0] n12138_o;
  wire [5:0] n12140_o;
  wire n12142_o;
  wire [5:0] n12143_o;
  wire n12144_o;
  wire [5:0] n12145_o;
  wire n12146_o;
  wire [31:0] n12147_o;
  wire [31:0] n12148_o;
  wire [31:0] n12149_o;
  localparam [32:0] n12150_o = 33'b000000000000000000000000000000000;
  wire n12151_o;
  wire n12153_o;
  wire n12154_o;
  wire n12155_o;
  wire n12156_o;
  wire n12157_o;
  wire [31:0] n12158_o;
  wire [31:0] n12159_o;
  wire n12160_o;
  wire n12162_o;
  wire n12164_o;
  wire [32:0] n12166_o;
  wire [1:0] n12167_o;
  wire n12168_o;
  localparam [23:0] n12169_o = 24'b000000000000000000000000;
  localparam [23:0] n12170_o = 24'b000000000000000000000000;
  wire n12172_o;
  wire n12173_o;
  wire n12174_o;
  wire n12175_o;
  wire [22:0] n12176_o;
  wire n12178_o;
  wire n12179_o;
  localparam [15:0] n12180_o = 16'b0000000000000000;
  wire n12183_o;
  wire n12184_o;
  wire n12185_o;
  wire n12186_o;
  wire [14:0] n12187_o;
  wire n12189_o;
  wire n12191_o;
  wire n12192_o;
  wire n12193_o;
  wire n12195_o;
  wire n12196_o;
  wire n12197_o;
  wire n12198_o;
  wire n12200_o;
  wire [2:0] n12201_o;
  wire n12202_o;
  reg n12203_o;
  wire [6:0] n12204_o;
  wire [6:0] n12205_o;
  reg [6:0] n12206_o;
  wire n12207_o;
  wire n12208_o;
  reg n12209_o;
  wire [14:0] n12210_o;
  wire [14:0] n12211_o;
  reg [14:0] n12212_o;
  wire n12213_o;
  reg n12214_o;
  wire [7:0] n12216_o;
  reg n12220_o;
  wire [7:0] n12221_o;
  wire [7:0] n12222_o;
  wire [7:0] n12223_o;
  wire [7:0] n12224_o;
  reg [7:0] n12225_o;
  wire [15:0] n12226_o;
  wire [15:0] n12227_o;
  wire [15:0] n12228_o;
  wire [15:0] n12229_o;
  reg [15:0] n12230_o;
  wire [7:0] n12234_o;
  wire [7:0] n12235_o;
  wire [7:0] n12236_o;
  wire [65:0] n12238_o;
  wire [30:0] n12239_o;
  wire [31:0] n12240_o;
  wire [65:0] n12241_o;
  wire n12245_o;
  wire [7:0] n12246_o;
  wire [7:0] n12247_o;
  wire n12248_o;
  wire [7:0] n12249_o;
  wire [7:0] n12250_o;
  wire n12251_o;
  wire [7:0] n12252_o;
  wire [7:0] n12253_o;
  wire [7:0] n12254_o;
  wire [7:0] n12255_o;
  wire [7:0] n12256_o;
  wire [7:0] n12257_o;
  wire n12258_o;
  wire n12259_o;
  wire n12260_o;
  wire n12261_o;
  wire [7:0] n12262_o;
  wire n12264_o;
  wire [7:0] n12266_o;
  wire n12268_o;
  wire [15:0] n12270_o;
  wire n12272_o;
  wire n12275_o;
  wire [1:0] n12276_o;
  wire [1:0] n12278_o;
  wire [2:0] n12279_o;
  wire [2:0] n12281_o;
  wire [2:0] n12283_o;
  wire n12286_o;
  wire n12287_o;
  wire n12288_o;
  wire [1:0] n12289_o;
  wire n12290_o;
  wire [2:0] n12291_o;
  wire n12292_o;
  wire [3:0] n12293_o;
  wire n12294_o;
  wire n12295_o;
  wire n12296_o;
  wire [1:0] n12297_o;
  wire [1:0] n12298_o;
  wire [1:0] n12299_o;
  wire [1:0] n12300_o;
  wire n12302_o;
  wire n12303_o;
  wire n12304_o;
  wire n12305_o;
  wire n12306_o;
  wire [1:0] n12307_o;
  wire n12308_o;
  wire [2:0] n12309_o;
  wire n12310_o;
  wire [3:0] n12311_o;
  wire n12312_o;
  wire n12313_o;
  wire [1:0] n12314_o;
  wire n12315_o;
  wire [2:0] n12316_o;
  wire n12317_o;
  wire [3:0] n12318_o;
  wire [3:0] n12319_o;
  wire [3:0] n12320_o;
  wire [3:0] n12321_o;
  wire n12323_o;
  wire n12324_o;
  wire n12327_o;
  wire n12330_o;
  wire n12331_o;
  wire n12332_o;
  wire n12333_o;
  wire n12334_o;
  wire n12335_o;
  wire n12337_o;
  wire n12338_o;
  wire n12340_o;
  wire n12341_o;
  wire n12342_o;
  wire n12343_o;
  wire n12344_o;
  wire [1:0] n12346_o;
  wire [3:0] n12348_o;
  wire [3:0] n12350_o;
  wire [3:0] n12351_o;
  wire [3:0] n12352_o;
  wire [3:0] n12353_o;
  wire [3:0] n12354_o;
  wire [3:0] n12355_o;
  wire [3:0] n12356_o;
  wire n12357_o;
  wire n12358_o;
  wire [3:0] n12359_o;
  wire n12360_o;
  wire n12361_o;
  wire n12362_o;
  wire n12364_o;
  wire n12365_o;
  wire n12366_o;
  wire n12367_o;
  wire n12368_o;
  wire n12369_o;
  wire n12370_o;
  wire n12371_o;
  wire n12372_o;
  wire n12373_o;
  wire n12374_o;
  wire n12375_o;
  wire n12376_o;
  wire n12377_o;
  wire n12378_o;
  wire n12379_o;
  wire n12380_o;
  wire n12381_o;
  wire n12383_o;
  wire n12385_o;
  wire n12387_o;
  wire n12388_o;
  wire n12389_o;
  wire [1:0] n12390_o;
  wire [3:0] n12392_o;
  wire n12393_o;
  wire n12394_o;
  wire [1:0] n12395_o;
  wire [3:0] n12397_o;
  wire [3:0] n12398_o;
  wire [3:0] n12399_o;
  wire n12400_o;
  wire n12402_o;
  wire n12403_o;
  wire n12404_o;
  wire n12405_o;
  wire n12406_o;
  wire n12409_o;
  wire n12411_o;
  wire n12412_o;
  wire n12413_o;
  wire n12415_o;
  wire n12416_o;
  wire n12417_o;
  wire n12418_o;
  wire n12419_o;
  wire n12420_o;
  wire n12421_o;
  wire n12422_o;
  wire n12423_o;
  wire n12424_o;
  wire n12425_o;
  wire n12426_o;
  wire n12427_o;
  wire n12428_o;
  wire n12430_o;
  wire n12431_o;
  wire n12434_o;
  wire n12435_o;
  wire n12436_o;
  wire n12437_o;
  wire n12438_o;
  wire [1:0] n12439_o;
  wire n12441_o;
  wire n12442_o;
  wire n12443_o;
  wire n12444_o;
  wire n12445_o;
  wire n12448_o;
  wire n12449_o;
  wire [1:0] n12450_o;
  wire n12451_o;
  wire n12452_o;
  wire n12453_o;
  wire n12454_o;
  wire n12455_o;
  wire n12456_o;
  wire n12457_o;
  wire n12458_o;
  wire n12459_o;
  wire n12460_o;
  wire n12461_o;
  wire n12462_o;
  wire n12463_o;
  wire n12464_o;
  wire n12465_o;
  wire n12466_o;
  wire n12467_o;
  wire n12468_o;
  wire n12469_o;
  wire n12470_o;
  wire n12471_o;
  wire n12472_o;
  wire n12474_o;
  wire n12475_o;
  wire n12476_o;
  wire n12477_o;
  wire n12478_o;
  wire n12479_o;
  wire n12481_o;
  wire n12482_o;
  wire n12483_o;
  wire n12484_o;
  wire [15:0] n12485_o;
  wire n12487_o;
  wire n12489_o;
  wire [15:0] n12490_o;
  wire n12492_o;
  wire n12493_o;
  wire n12494_o;
  wire n12497_o;
  wire [3:0] n12500_o;
  wire [3:0] n12501_o;
  wire [3:0] n12502_o;
  wire [3:0] n12503_o;
  wire [3:0] n12504_o;
  wire [3:0] n12505_o;
  wire [3:0] n12506_o;
  wire [3:0] n12507_o;
  wire [3:0] n12508_o;
  wire [1:0] n12509_o;
  wire [1:0] n12510_o;
  wire [1:0] n12511_o;
  wire [1:0] n12512_o;
  wire [1:0] n12513_o;
  wire [1:0] n12514_o;
  wire [1:0] n12515_o;
  wire n12516_o;
  wire n12517_o;
  wire n12518_o;
  wire n12519_o;
  wire n12520_o;
  wire n12521_o;
  wire n12522_o;
  wire n12523_o;
  wire n12524_o;
  wire [3:0] n12525_o;
  wire [3:0] n12526_o;
  wire [3:0] n12527_o;
  wire [3:0] n12528_o;
  wire [3:0] n12529_o;
  wire [3:0] n12530_o;
  wire [3:0] n12531_o;
  wire [3:0] n12532_o;
  wire [3:0] n12533_o;
  wire [3:0] n12534_o;
  wire [3:0] n12535_o;
  wire [3:0] n12536_o;
  wire [3:0] n12537_o;
  wire [4:0] n12538_o;
  wire [4:0] n12539_o;
  wire [4:0] n12540_o;
  wire [4:0] n12541_o;
  wire [4:0] n12542_o;
  wire [4:0] n12543_o;
  wire [4:0] n12544_o;
  wire [3:0] n12545_o;
  wire [3:0] n12546_o;
  wire [3:0] n12547_o;
  wire n12548_o;
  wire n12549_o;
  wire n12550_o;
  wire n12551_o;
  wire n12552_o;
  wire n12553_o;
  wire n12554_o;
  wire [3:0] n12555_o;
  wire [4:0] n12556_o;
  wire [4:0] n12557_o;
  wire [4:0] n12558_o;
  wire [2:0] n12559_o;
  wire [2:0] n12560_o;
  wire [2:0] n12561_o;
  wire [2:0] n12562_o;
  wire [2:0] n12563_o;
  wire [2:0] n12564_o;
  wire [2:0] n12565_o;
  wire [3:0] n12571_o;
  wire [7:0] n12572_o;
  wire [3:0] n12574_o;
  wire n12575_o;
  localparam [7:0] n12576_o = 8'b00000000;
  wire [3:0] n12578_o;
  wire n12579_o;
  wire [4:0] n12581_o;
  wire [4:0] n12582_o;
  wire [4:0] n12583_o;
  wire [4:0] n12584_o;
  wire [4:0] n12585_o;
  wire [7:0] n12586_o;
  wire n12593_o;
  wire n12594_o;
  wire n12595_o;
  wire [31:0] n12598_o;
  wire n12599_o;
  wire n12600_o;
  wire [31:0] n12603_o;
  wire [15:0] n12604_o;
  wire [15:0] n12605_o;
  wire n12606_o;
  wire n12607_o;
  wire [15:0] n12610_o;
  wire n12611_o;
  wire n12612_o;
  wire [15:0] n12615_o;
  wire [31:0] n12616_o;
  wire [31:0] n12617_o;
  wire [31:0] n12618_o;
  wire [31:0] n12619_o;
  wire [15:0] n12620_o;
  wire [47:0] n12621_o;
  wire [15:0] n12622_o;
  wire [63:0] n12623_o;
  wire [15:0] n12624_o;
  wire [47:0] n12625_o;
  wire [15:0] n12626_o;
  wire [63:0] n12627_o;
  wire [127:0] n12628_o;
  wire [127:0] n12629_o;
  wire [127:0] n12630_o;
  wire [31:0] n12631_o;
  wire n12633_o;
  wire n12634_o;
  wire n12635_o;
  wire n12636_o;
  wire n12637_o;
  wire n12638_o;
  wire [31:0] n12639_o;
  wire n12641_o;
  wire n12642_o;
  wire n12643_o;
  wire n12644_o;
  wire n12645_o;
  wire n12648_o;
  wire [31:0] n12653_o;
  wire n12661_o;
  wire n12662_o;
  wire n12663_o;
  wire n12664_o;
  wire n12665_o;
  wire n12666_o;
  wire n12667_o;
  wire n12668_o;
  wire n12670_o;
  wire n12671_o;
  wire n12672_o;
  wire n12673_o;
  wire n12674_o;
  wire n12675_o;
  wire n12676_o;
  wire n12677_o;
  wire n12678_o;
  wire n12679_o;
  wire n12680_o;
  wire n12681_o;
  wire n12682_o;
  wire n12683_o;
  wire n12684_o;
  wire n12685_o;
  wire n12686_o;
  wire n12687_o;
  wire n12688_o;
  wire n12689_o;
  wire n12690_o;
  wire n12691_o;
  wire n12692_o;
  wire n12693_o;
  wire n12694_o;
  wire n12695_o;
  wire n12696_o;
  wire n12697_o;
  wire n12698_o;
  wire n12699_o;
  wire n12700_o;
  wire n12701_o;
  wire n12702_o;
  wire n12703_o;
  wire n12704_o;
  wire n12705_o;
  wire n12706_o;
  wire n12707_o;
  wire n12708_o;
  wire n12709_o;
  wire n12710_o;
  wire n12711_o;
  wire n12712_o;
  wire n12713_o;
  wire n12714_o;
  wire n12715_o;
  wire n12716_o;
  wire n12717_o;
  wire n12718_o;
  wire n12719_o;
  wire n12720_o;
  wire n12721_o;
  wire n12722_o;
  wire n12723_o;
  wire n12724_o;
  wire n12725_o;
  wire n12726_o;
  wire n12727_o;
  wire n12728_o;
  wire n12729_o;
  wire n12730_o;
  wire n12731_o;
  wire n12732_o;
  wire n12733_o;
  wire [3:0] n12734_o;
  wire [3:0] n12735_o;
  wire [3:0] n12736_o;
  wire [3:0] n12737_o;
  wire [3:0] n12738_o;
  wire [3:0] n12739_o;
  wire [3:0] n12740_o;
  wire [3:0] n12741_o;
  wire [15:0] n12742_o;
  wire [15:0] n12743_o;
  wire [31:0] n12744_o;
  wire n12745_o;
  wire n12747_o;
  wire n12748_o;
  wire n12749_o;
  wire n12750_o;
  wire n12751_o;
  wire [31:0] n12752_o;
  wire n12753_o;
  wire n12754_o;
  wire [63:0] n12755_o;
  wire [15:0] n12756_o;
  wire [15:0] n12757_o;
  wire [31:0] n12758_o;
  wire [31:0] n12759_o;
  wire [15:0] n12760_o;
  wire [15:0] n12761_o;
  wire [15:0] n12762_o;
  wire n12764_o;
  wire n12765_o;
  wire n12766_o;
  wire [15:0] n12767_o;
  wire [15:0] n12769_o;
  wire n12770_o;
  wire n12771_o;
  wire [32:0] n12772_o;
  wire [32:0] n12774_o;
  wire [32:0] n12775_o;
  wire [32:0] n12776_o;
  wire [16:0] n12778_o;
  wire [15:0] n12779_o;
  wire [32:0] n12780_o;
  wire [32:0] n12781_o;
  wire [32:0] n12782_o;
  wire n12783_o;
  wire [31:0] n12784_o;
  wire [31:0] n12785_o;
  wire [31:0] n12786_o;
  wire [30:0] n12787_o;
  wire n12788_o;
  wire [31:0] n12789_o;
  wire [31:0] n12790_o;
  wire [31:0] n12792_o;
  wire [31:0] n12793_o;
  wire [31:0] n12794_o;
  wire n12795_o;
  wire n12796_o;
  wire n12797_o;
  wire n12798_o;
  wire n12799_o;
  wire n12800_o;
  wire n12801_o;
  wire n12802_o;
  wire n12803_o;
  wire n12804_o;
  wire n12805_o;
  wire n12806_o;
  wire n12808_o;
  wire n12811_o;
  wire n12817_o;
  wire n12820_o;
  wire n12821_o;
  wire n12822_o;
  wire [63:0] n12824_o;
  wire [63:0] n12825_o;
  wire n12828_o;
  wire n12829_o;
  wire n12830_o;
  wire [63:0] n12831_o;
  wire n12833_o;
  wire n12836_o;
  wire n12837_o;
  wire n12838_o;
  wire n12839_o;
  wire [31:0] n12840_o;
  wire [32:0] n12842_o;
  wire [16:0] n12844_o;
  wire [15:0] n12845_o;
  wire [32:0] n12846_o;
  wire [32:0] n12847_o;
  wire n12850_o;
  wire n12851_o;
  wire [31:0] n12852_o;
  wire [31:0] n12854_o;
  wire [31:0] n12855_o;
  wire [31:0] n12856_o;
  wire [63:0] n12857_o;
  wire n12859_o;
  wire n12860_o;
  wire n12862_o;
  wire n12863_o;
  wire n12866_o;
  wire [31:0] n12876_o;
  wire [2:0] n12877_o;
  wire [3:0] n12878_o;
  reg [3:0] n12879_q;
  wire [8:0] n12880_o;
  wire [63:0] n12881_o;
  reg [63:0] n12882_q;
  wire n12883_o;
  reg n12884_q;
  reg n12885_q;
  wire n12887_o;
  reg n12888_q;
  wire n12889_o;
  reg n12890_q;
  wire [31:0] n12894_o;
  wire [31:0] n12895_o;
  reg [31:0] n12896_q;
  wire [63:0] n12898_o;
  wire [63:0] n12900_o;
  reg [63:0] n12901_q;
  wire [63:0] n12902_o;
  wire n12904_o;
  reg n12905_q;
  wire [32:0] n12906_o;
  reg [32:0] n12907_q;
  wire n12908_o;
  reg n12909_q;
  wire [63:0] n12910_o;
  wire n12911_o;
  reg n12912_q;
  wire n12913_o;
  reg n12914_q;
  wire [31:0] n12917_o;
  wire [39:0] n12919_o;
  wire [31:0] n12920_o;
  wire [39:0] n12922_o;
  wire [4:0] n12923_o;
  wire n12924_o;
  reg n12925_q;
  wire n12926_o;
  reg n12927_q;
  wire n12928_o;
  reg n12929_q;
  wire n12930_o;
  reg n12931_q;
  wire n12932_o;
  reg n12933_q;
  wire n12934_o;
  reg n12935_q;
  wire n12936_o;
  reg n12937_q;
  wire [32:0] n12939_o;
  wire [32:0] n12940_o;
  wire [32:0] n12941_o;
  wire [31:0] n12942_o;
  wire [7:0] n12943_o;
  reg [7:0] n12944_q;
  reg [7:0] n12945_q;
  wire n12946_o;
  wire n12947_o;
  wire n12948_o;
  wire n12949_o;
  wire n12950_o;
  wire n12951_o;
  wire n12952_o;
  wire n12953_o;
  wire n12954_o;
  wire n12955_o;
  wire n12956_o;
  wire n12957_o;
  wire n12958_o;
  wire n12959_o;
  wire n12960_o;
  wire n12961_o;
  wire n12962_o;
  wire n12963_o;
  wire n12964_o;
  wire n12965_o;
  wire n12966_o;
  wire n12967_o;
  wire n12968_o;
  wire n12969_o;
  wire n12970_o;
  wire n12971_o;
  wire n12972_o;
  wire n12973_o;
  wire n12974_o;
  wire n12975_o;
  wire n12976_o;
  wire n12977_o;
  wire [1:0] n12978_o;
  reg n12979_o;
  wire [1:0] n12980_o;
  reg n12981_o;
  wire [1:0] n12982_o;
  reg n12983_o;
  wire [1:0] n12984_o;
  reg n12985_o;
  wire [1:0] n12986_o;
  reg n12987_o;
  wire [1:0] n12988_o;
  reg n12989_o;
  wire [1:0] n12990_o;
  reg n12991_o;
  wire [1:0] n12992_o;
  reg n12993_o;
  wire [1:0] n12994_o;
  reg n12995_o;
  wire [1:0] n12996_o;
  reg n12997_o;
  wire n12998_o;
  wire n12999_o;
  wire n13000_o;
  wire n13001_o;
  wire n13002_o;
  wire n13003_o;
  wire n13004_o;
  wire n13005_o;
  wire n13006_o;
  wire n13007_o;
  wire n13008_o;
  wire n13009_o;
  wire n13010_o;
  wire n13011_o;
  wire n13012_o;
  wire n13013_o;
  wire n13014_o;
  wire n13015_o;
  wire n13016_o;
  wire n13017_o;
  wire n13018_o;
  wire n13019_o;
  wire n13020_o;
  wire n13021_o;
  wire n13022_o;
  wire n13023_o;
  wire n13024_o;
  wire n13025_o;
  wire n13026_o;
  wire n13027_o;
  wire n13028_o;
  wire n13029_o;
  wire n13030_o;
  wire n13031_o;
  wire n13032_o;
  wire n13033_o;
  wire n13034_o;
  wire n13035_o;
  wire n13036_o;
  wire n13037_o;
  wire n13038_o;
  wire n13039_o;
  wire n13040_o;
  wire n13041_o;
  wire n13042_o;
  wire n13043_o;
  wire n13044_o;
  wire n13045_o;
  wire n13046_o;
  wire n13047_o;
  wire n13048_o;
  wire n13049_o;
  wire n13050_o;
  wire n13051_o;
  wire n13052_o;
  wire n13053_o;
  wire n13054_o;
  wire n13055_o;
  wire n13056_o;
  wire n13057_o;
  wire n13058_o;
  wire n13059_o;
  wire n13060_o;
  wire n13061_o;
  wire n13062_o;
  wire n13063_o;
  wire n13064_o;
  wire n13065_o;
  wire n13066_o;
  wire n13067_o;
  wire n13068_o;
  wire n13069_o;
  wire n13070_o;
  wire n13071_o;
  wire n13072_o;
  wire n13073_o;
  wire n13074_o;
  wire n13075_o;
  wire n13076_o;
  wire n13077_o;
  wire n13078_o;
  wire n13079_o;
  wire n13080_o;
  wire n13081_o;
  wire n13082_o;
  wire n13083_o;
  wire n13084_o;
  wire n13085_o;
  wire n13086_o;
  wire n13087_o;
  wire n13088_o;
  wire n13089_o;
  wire n13090_o;
  wire n13091_o;
  wire n13092_o;
  wire n13093_o;
  wire n13094_o;
  wire n13095_o;
  wire n13096_o;
  wire n13097_o;
  wire n13098_o;
  wire n13099_o;
  wire n13100_o;
  wire n13101_o;
  wire n13102_o;
  wire n13103_o;
  wire n13104_o;
  wire n13105_o;
  wire n13106_o;
  wire n13107_o;
  wire n13108_o;
  wire n13109_o;
  wire n13110_o;
  wire n13111_o;
  wire n13112_o;
  wire n13113_o;
  wire n13114_o;
  wire n13115_o;
  wire n13116_o;
  wire n13117_o;
  wire n13118_o;
  wire n13119_o;
  wire n13120_o;
  wire n13121_o;
  wire n13122_o;
  wire n13123_o;
  wire n13124_o;
  wire n13125_o;
  wire n13126_o;
  wire n13127_o;
  wire n13128_o;
  wire n13129_o;
  wire n13130_o;
  wire n13131_o;
  wire n13132_o;
  wire n13133_o;
  wire [31:0] n13134_o;
  wire n13135_o;
  wire n13136_o;
  wire n13137_o;
  wire n13138_o;
  wire n13139_o;
  wire n13140_o;
  wire n13141_o;
  wire n13142_o;
  wire n13143_o;
  wire n13144_o;
  wire n13145_o;
  wire n13146_o;
  wire n13147_o;
  wire n13148_o;
  wire n13149_o;
  wire n13150_o;
  wire n13151_o;
  wire n13152_o;
  wire n13153_o;
  wire n13154_o;
  wire n13155_o;
  wire n13156_o;
  wire n13157_o;
  wire n13158_o;
  wire n13159_o;
  wire n13160_o;
  wire n13161_o;
  wire n13162_o;
  wire n13163_o;
  wire n13164_o;
  wire n13165_o;
  wire n13166_o;
  wire [1:0] n13167_o;
  reg n13168_o;
  wire [1:0] n13169_o;
  reg n13170_o;
  wire [1:0] n13171_o;
  reg n13172_o;
  wire [1:0] n13173_o;
  reg n13174_o;
  wire [1:0] n13175_o;
  reg n13176_o;
  wire [1:0] n13177_o;
  reg n13178_o;
  wire [1:0] n13179_o;
  reg n13180_o;
  wire [1:0] n13181_o;
  reg n13182_o;
  wire [1:0] n13183_o;
  reg n13184_o;
  wire [1:0] n13185_o;
  reg n13186_o;
  wire n13187_o;
  wire n13188_o;
  wire n13189_o;
  wire n13190_o;
  wire n13191_o;
  wire n13192_o;
  wire n13193_o;
  wire n13194_o;
  wire n13195_o;
  wire n13196_o;
  wire n13197_o;
  wire n13198_o;
  wire n13199_o;
  wire n13200_o;
  wire n13201_o;
  wire n13202_o;
  wire n13203_o;
  wire n13204_o;
  wire n13205_o;
  wire n13206_o;
  wire n13207_o;
  wire n13208_o;
  wire n13209_o;
  wire n13210_o;
  wire n13211_o;
  wire n13212_o;
  wire n13213_o;
  wire n13214_o;
  wire n13215_o;
  wire n13216_o;
  wire n13217_o;
  wire n13218_o;
  wire n13219_o;
  wire n13220_o;
  wire n13221_o;
  wire n13222_o;
  wire n13223_o;
  wire n13224_o;
  wire n13225_o;
  wire n13226_o;
  wire n13227_o;
  wire n13228_o;
  wire n13229_o;
  wire n13230_o;
  wire n13231_o;
  wire n13232_o;
  wire n13233_o;
  wire n13234_o;
  wire n13235_o;
  wire n13236_o;
  wire n13237_o;
  wire n13238_o;
  wire n13239_o;
  wire n13240_o;
  wire n13241_o;
  wire n13242_o;
  wire n13243_o;
  wire n13244_o;
  wire n13245_o;
  wire n13246_o;
  wire n13247_o;
  wire n13248_o;
  wire n13249_o;
  wire n13250_o;
  wire n13251_o;
  wire n13252_o;
  wire n13253_o;
  wire n13254_o;
  wire n13255_o;
  wire n13256_o;
  wire n13257_o;
  wire n13258_o;
  wire n13259_o;
  wire n13260_o;
  wire n13261_o;
  wire n13262_o;
  wire n13263_o;
  wire n13264_o;
  wire n13265_o;
  wire n13266_o;
  wire n13267_o;
  wire n13268_o;
  wire n13269_o;
  wire n13270_o;
  wire n13271_o;
  wire n13272_o;
  wire n13273_o;
  wire n13274_o;
  wire n13275_o;
  wire n13276_o;
  wire n13277_o;
  wire n13278_o;
  wire n13279_o;
  wire n13280_o;
  wire n13281_o;
  wire n13282_o;
  wire n13283_o;
  wire n13284_o;
  wire n13285_o;
  wire n13286_o;
  wire n13287_o;
  wire n13288_o;
  wire n13289_o;
  wire n13290_o;
  wire n13291_o;
  wire n13292_o;
  wire n13293_o;
  wire n13294_o;
  wire n13295_o;
  wire n13296_o;
  wire n13297_o;
  wire n13298_o;
  wire n13299_o;
  wire n13300_o;
  wire n13301_o;
  wire n13302_o;
  wire n13303_o;
  wire n13304_o;
  wire n13305_o;
  wire n13306_o;
  wire n13307_o;
  wire n13308_o;
  wire n13309_o;
  wire n13310_o;
  wire n13311_o;
  wire n13312_o;
  wire n13313_o;
  wire n13314_o;
  wire n13315_o;
  wire n13316_o;
  wire n13317_o;
  wire n13318_o;
  wire n13319_o;
  wire n13320_o;
  wire n13321_o;
  wire n13322_o;
  wire n13323_o;
  wire n13324_o;
  wire n13325_o;
  wire n13326_o;
  wire n13327_o;
  wire n13328_o;
  wire n13329_o;
  wire n13330_o;
  wire n13331_o;
  wire n13332_o;
  wire n13333_o;
  wire n13334_o;
  wire n13335_o;
  wire n13336_o;
  wire [33:0] n13337_o;
  assign bf_ext_out = n12944_q;
  assign set_v_flag = n12811_o;
  assign flags = n12945_q;
  assign c_out = n10188_o;
  assign addsub_q = n10166_o;
  assign aluout = n9948_o;
  /* TG68K_ALU.vhd:86:16  */
  assign op1in = n12876_o; // (signal)
  /* TG68K_ALU.vhd:87:16  */
  assign addsub_a = n10054_o; // (signal)
  /* TG68K_ALU.vhd:88:16  */
  assign addsub_b = n10137_o; // (signal)
  /* TG68K_ALU.vhd:89:16  */
  assign notaddsub_b = n10149_o; // (signal)
  /* TG68K_ALU.vhd:90:16  */
  assign add_result = n10154_o; // (signal)
  /* TG68K_ALU.vhd:91:16  */
  assign addsub_ofl = n12877_o; // (signal)
  /* TG68K_ALU.vhd:92:16  */
  assign opaddsub = n10116_o; // (signal)
  /* TG68K_ALU.vhd:93:16  */
  assign c_in = n12878_o; // (signal)
  /* TG68K_ALU.vhd:94:16  */
  assign flag_z = n12283_o; // (signal)
  /* TG68K_ALU.vhd:95:16  */
  assign set_flags = n12321_o; // (signal)
  /* TG68K_ALU.vhd:96:16  */
  assign ccrin = n12257_o; // (signal)
  /* TG68K_ALU.vhd:97:16  */
  assign last_flags1 = n12879_q; // (signal)
  /* TG68K_ALU.vhd:100:16  */
  assign bcd_pur = n10194_o; // (signal)
  /* TG68K_ALU.vhd:101:16  */
  assign bcd_kor = n12880_o; // (signal)
  /* TG68K_ALU.vhd:102:16  */
  assign halve_carry = n10199_o; // (signal)
  /* TG68K_ALU.vhd:103:16  */
  assign vflag_a = n10252_o; // (signal)
  /* TG68K_ALU.vhd:104:16  */
  assign bcd_a_carry = n10255_o; // (signal)
  /* TG68K_ALU.vhd:105:16  */
  assign bcd_a = n10249_o; // (signal)
  /* TG68K_ALU.vhd:106:16  */
  assign result_mulu = n12630_o; // (signal)
  /* TG68K_ALU.vhd:107:16  */
  assign result_div = n12882_q; // (signal)
  /* TG68K_ALU.vhd:108:16  */
  assign result_div_pre = n12794_o; // (signal)
  /* TG68K_ALU.vhd:109:16  */
  assign set_mv_flag = n12648_o; // (signal)
  /* TG68K_ALU.vhd:110:16  */
  assign v_flag = n12884_q; // (signal)
  /* TG68K_ALU.vhd:112:16  */
  assign rot_rot = n11745_o; // (signal)
  /* TG68K_ALU.vhd:115:16  */
  assign rot_x = n11798_o; // (signal)
  /* TG68K_ALU.vhd:116:16  */
  assign rot_c = n11799_o; // (signal)
  /* TG68K_ALU.vhd:117:16  */
  assign rot_out = n11800_o; // (signal)
  /* TG68K_ALU.vhd:118:16  */
  assign asl_vflag = n12885_q; // (signal)
  /* TG68K_ALU.vhd:120:16  */
  assign bit_number = n10296_o; // (signal)
  /* TG68K_ALU.vhd:121:16  */
  assign bits_out = n13134_o; // (signal)
  /* TG68K_ALU.vhd:122:16  */
  assign one_bit_in = n12999_o; // (signal)
  /* TG68K_ALU.vhd:123:16  */
  assign bchg = n12888_q; // (signal)
  /* TG68K_ALU.vhd:124:16  */
  assign bset = n12890_q; // (signal)
  /* TG68K_ALU.vhd:129:16  */
  assign mulu_reg = n12898_o; // (signal)
  /* TG68K_ALU.vhd:131:16  */
  assign faktora = n12617_o; // (signal)
  /* TG68K_ALU.vhd:132:16  */
  assign faktorb = n12619_o; // (signal)
  /* TG68K_ALU.vhd:134:16  */
  assign div_reg = n12901_q; // (signal)
  /* TG68K_ALU.vhd:135:16  */
  assign div_quot = n12902_o; // (signal)
  /* TG68K_ALU.vhd:137:16  */
  assign div_neg = n12905_q; // (signal)
  /* TG68K_ALU.vhd:138:16  */
  assign div_bit = n12783_o; // (signal)
  /* TG68K_ALU.vhd:139:16  */
  assign div_sub = n12782_o; // (signal)
  /* TG68K_ALU.vhd:140:16  */
  assign div_over = n12907_q; // (signal)
  /* TG68K_ALU.vhd:141:16  */
  assign nozero = n12909_q; // (signal)
  /* TG68K_ALU.vhd:142:16  */
  assign div_qsign = n12754_o; // (signal)
  /* TG68K_ALU.vhd:143:16  */
  assign dividend = n12910_o; // (signal)
  /* TG68K_ALU.vhd:144:16  */
  assign divs = n12668_o; // (signal)
  /* TG68K_ALU.vhd:145:16  */
  assign signedop = n12912_q; // (signal)
  /* TG68K_ALU.vhd:146:16  */
  assign op1_sign = n12914_q; // (signal)
  /* TG68K_ALU.vhd:148:16  */
  assign op2outext = n12769_o; // (signal)
  /* TG68K_ALU.vhd:151:16  */
  assign datareg = n12917_o; // (signal)
  /* TG68K_ALU.vhd:153:16  */
  assign bf_datareg = n10855_o; // (signal)
  /* TG68K_ALU.vhd:154:16  */
  assign result = n12919_o; // (signal)
  /* TG68K_ALU.vhd:155:16  */
  assign result_tmp = n10944_o; // (signal)
  /* TG68K_ALU.vhd:156:16  */
  assign unshifted_bitmask = n12920_o; // (signal)
  /* TG68K_ALU.vhd:158:16  */
  assign inmux0 = n10910_o; // (signal)
  /* TG68K_ALU.vhd:159:16  */
  assign inmux1 = n10915_o; // (signal)
  /* TG68K_ALU.vhd:160:16  */
  assign inmux2 = n10920_o; // (signal)
  /* TG68K_ALU.vhd:161:16  */
  assign inmux3 = n10926_o; // (signal)
  /* TG68K_ALU.vhd:162:16  */
  assign shifted_bitmask = n10900_o; // (signal)
  /* TG68K_ALU.vhd:163:16  */
  assign bitmaskmux0 = n10887_o; // (signal)
  /* TG68K_ALU.vhd:164:16  */
  assign bitmaskmux1 = n10876_o; // (signal)
  /* TG68K_ALU.vhd:165:16  */
  assign bitmaskmux2 = n10865_o; // (signal)
  /* TG68K_ALU.vhd:166:16  */
  assign bitmaskmux3 = n10860_o; // (signal)
  /* TG68K_ALU.vhd:167:16  */
  assign bf_set2 = n10931_o; // (signal)
  /* TG68K_ALU.vhd:168:16  */
  assign shift = n12922_o; // (signal)
  /* TG68K_ALU.vhd:169:16  */
  assign bf_firstbit = n11614_o; // (signal)
  /* TG68K_ALU.vhd:170:16  */
  assign mux = n11691_o; // (signal)
  /* TG68K_ALU.vhd:171:16  */
  assign bitnr = n12923_o; // (signal)
  /* TG68K_ALU.vhd:172:16  */
  assign mask = datareg; // (signal)
  /* TG68K_ALU.vhd:173:16  */
  assign mask_not_zero = n11726_o; // (signal)
  /* TG68K_ALU.vhd:174:16  */
  assign bf_bset = n12925_q; // (signal)
  /* TG68K_ALU.vhd:175:16  */
  assign bf_nflag = n13188_o; // (signal)
  /* TG68K_ALU.vhd:176:16  */
  assign bf_bchg = n12927_q; // (signal)
  /* TG68K_ALU.vhd:177:16  */
  assign bf_ins = n12929_q; // (signal)
  /* TG68K_ALU.vhd:178:16  */
  assign bf_exts = n12931_q; // (signal)
  /* TG68K_ALU.vhd:179:16  */
  assign bf_fffo = n12933_q; // (signal)
  /* TG68K_ALU.vhd:180:16  */
  assign bf_d32 = n12935_q; // (signal)
  /* TG68K_ALU.vhd:181:16  */
  assign bf_s32 = n12937_q; // (signal)
  /* TG68K_ALU.vhd:187:16  */
  assign hot_msb = n13337_o; // (signal)
  /* TG68K_ALU.vhd:188:16  */
  assign vector = n12939_o; // (signal)
  /* TG68K_ALU.vhd:189:16  */
  assign result_bs = n12241_o; // (signal)
  /* TG68K_ALU.vhd:190:16  */
  assign bit_nr = n12145_o; // (signal)
  /* TG68K_ALU.vhd:191:16  */
  assign bit_msb = n11868_o; // (signal)
  /* TG68K_ALU.vhd:192:16  */
  assign bs_shift = n11858_o; // (signal)
  /* TG68K_ALU.vhd:193:16  */
  assign bs_shift_mod = n12115_o; // (signal)
  /* TG68K_ALU.vhd:194:16  */
  assign asl_over = n11900_o; // (signal)
  /* TG68K_ALU.vhd:195:16  */
  assign asl_over_xor = n12940_o; // (signal)
  /* TG68K_ALU.vhd:196:16  */
  assign asr_sign = n12941_o; // (signal)
  /* TG68K_ALU.vhd:197:16  */
  assign msb = n12220_o; // (signal)
  /* TG68K_ALU.vhd:198:16  */
  assign ring = n11838_o; // (signal)
  /* TG68K_ALU.vhd:199:16  */
  assign alu = n12022_o; // (signal)
  /* TG68K_ALU.vhd:200:16  */
  assign bsout = n12942_o; // (signal)
  /* TG68K_ALU.vhd:201:16  */
  assign bs_v = n12035_o; // (signal)
  /* TG68K_ALU.vhd:202:16  */
  assign bs_c = n12162_o; // (signal)
  /* TG68K_ALU.vhd:203:16  */
  assign bs_x = n12037_o; // (signal)
  /* TG68K_ALU.vhd:215:35  */
  assign n9938_o = op1in[7];
  /* TG68K_ALU.vhd:215:39  */
  assign n9939_o = n9938_o | exec_tas;
  assign n9940_o = op1in[31:8];
  assign n9941_o = op1in[6:0];
  /* TG68K_ALU.vhd:216:24  */
  assign n9942_o = exec[76];
  /* TG68K_ALU.vhd:217:41  */
  assign n9943_o = result[31:0];
  /* TG68K_ALU.vhd:219:57  */
  assign n9944_o = {26'b0, bf_firstbit};  //  uext
  /* TG68K_ALU.vhd:219:57  */
  assign n9945_o = bf_ffo_offset - n9944_o;
  /* TG68K_ALU.vhd:218:25  */
  assign n9946_o = bf_fffo ? n9945_o : n9943_o;
  assign n9947_o = {n9940_o, n9939_o, n9941_o};
  /* TG68K_ALU.vhd:216:17  */
  assign n9948_o = n9942_o ? n9946_o : n9947_o;
  /* TG68K_ALU.vhd:224:24  */
  assign n9949_o = exec[12];
  /* TG68K_ALU.vhd:224:45  */
  assign n9950_o = exec[13];
  /* TG68K_ALU.vhd:224:38  */
  assign n9951_o = n9949_o | n9950_o;
  /* TG68K_ALU.vhd:225:51  */
  assign n9952_o = bcd_a[7:0];
  /* TG68K_ALU.vhd:226:27  */
  assign n9953_o = exec[20];
  /* TG68K_ALU.vhd:226:41  */
  assign n9955_o = 1'b1 & n9953_o;
  /* TG68K_ALU.vhd:234:40  */
  assign n9956_o = exec[67];
  /* TG68K_ALU.vhd:235:61  */
  assign n9957_o = result_mulu[31:0];
  /* TG68K_ALU.vhd:238:58  */
  assign n9958_o = mulu_reg[31:0];
  /* TG68K_ALU.vhd:234:33  */
  assign n9959_o = n9956_o ? n9957_o : n9958_o;
  /* TG68K_ALU.vhd:241:27  */
  assign n9960_o = exec[21];
  /* TG68K_ALU.vhd:241:41  */
  assign n9962_o = 1'b1 & n9960_o;
  /* TG68K_ALU.vhd:242:38  */
  assign n9963_o = exe_opcode[15];
  /* TG68K_ALU.vhd:242:47  */
  assign n9965_o = n9963_o | 1'b0;
  /* TG68K_ALU.vhd:244:52  */
  assign n9966_o = result_div[47:32];
  /* TG68K_ALU.vhd:244:77  */
  assign n9967_o = result_div[15:0];
  /* TG68K_ALU.vhd:244:66  */
  assign n9968_o = {n9966_o, n9967_o};
  /* TG68K_ALU.vhd:246:40  */
  assign n9969_o = exec[68];
  /* TG68K_ALU.vhd:247:60  */
  assign n9970_o = result_div[63:32];
  /* TG68K_ALU.vhd:249:60  */
  assign n9971_o = result_div[31:0];
  /* TG68K_ALU.vhd:246:33  */
  assign n9972_o = n9969_o ? n9970_o : n9971_o;
  /* TG68K_ALU.vhd:242:25  */
  assign n9973_o = n9965_o ? n9968_o : n9972_o;
  /* TG68K_ALU.vhd:252:27  */
  assign n9974_o = exec[5];
  /* TG68K_ALU.vhd:253:41  */
  assign n9975_o = op2out | op1out;
  /* TG68K_ALU.vhd:254:27  */
  assign n9976_o = exec[6];
  /* TG68K_ALU.vhd:255:41  */
  assign n9977_o = op2out & op1out;
  /* TG68K_ALU.vhd:256:27  */
  assign n9978_o = exec[16];
  assign n9979_o = {exe_condition, exe_condition, exe_condition, exe_condition};
  assign n9980_o = {exe_condition, exe_condition, exe_condition, exe_condition};
  assign n9981_o = {n9979_o, n9980_o};
  /* TG68K_ALU.vhd:258:27  */
  assign n9982_o = exec[7];
  /* TG68K_ALU.vhd:259:41  */
  assign n9983_o = op2out ^ op1out;
  /* TG68K_ALU.vhd:261:27  */
  assign n9984_o = exec[85];
  /* TG68K_ALU.vhd:264:27  */
  assign n9985_o = exec[9];
  /* TG68K_ALU.vhd:266:27  */
  assign n9986_o = exec[81];
  /* TG68K_ALU.vhd:268:27  */
  assign n9987_o = exec[15];
  /* TG68K_ALU.vhd:269:40  */
  assign n9988_o = op1out[15:0];
  /* TG68K_ALU.vhd:269:61  */
  assign n9989_o = op1out[31:16];
  /* TG68K_ALU.vhd:269:53  */
  assign n9990_o = {n9988_o, n9989_o};
  /* TG68K_ALU.vhd:270:27  */
  assign n9991_o = exec[14];
  /* TG68K_ALU.vhd:272:27  */
  assign n9992_o = exec[75];
  /* TG68K_ALU.vhd:274:27  */
  assign n9993_o = exec[2];
  /* TG68K_ALU.vhd:276:38  */
  assign n9994_o = exe_opcode[9];
  /* TG68K_ALU.vhd:276:25  */
  assign n9996_o = n9994_o ? 8'b00000000 : flagssr;
  /* TG68K_ALU.vhd:281:27  */
  assign n9997_o = exec[77];
  /* TG68K_ALU.vhd:282:54  */
  assign n9998_o = n10166_o[11:8];
  /* TG68K_ALU.vhd:282:78  */
  assign n9999_o = n10166_o[3:0];
  /* TG68K_ALU.vhd:282:68  */
  assign n10000_o = {n9998_o, n9999_o};
  assign n10001_o = n10166_o[7:0];
  /* TG68K_ALU.vhd:281:17  */
  assign n10002_o = n9997_o ? n10000_o : n10001_o;
  assign n10003_o = {n9996_o, n12945_q};
  assign n10004_o = n10003_o[7:0];
  /* TG68K_ALU.vhd:274:17  */
  assign n10005_o = n9993_o ? n10004_o : n10002_o;
  assign n10006_o = n10003_o[15:8];
  assign n10007_o = n10166_o[15:8];
  /* TG68K_ALU.vhd:274:17  */
  assign n10008_o = n9993_o ? n10006_o : n10007_o;
  assign n10009_o = {n10008_o, n10005_o};
  assign n10010_o = bf_datareg[15:0];
  /* TG68K_ALU.vhd:272:17  */
  assign n10011_o = n9992_o ? n10010_o : n10009_o;
  assign n10012_o = bf_datareg[31:16];
  assign n10013_o = n10166_o[31:16];
  /* TG68K_ALU.vhd:272:17  */
  assign n10014_o = n9992_o ? n10012_o : n10013_o;
  assign n10015_o = {n10014_o, n10011_o};
  /* TG68K_ALU.vhd:270:17  */
  assign n10016_o = n9991_o ? bits_out : n10015_o;
  /* TG68K_ALU.vhd:268:17  */
  assign n10017_o = n9987_o ? n9990_o : n10016_o;
  /* TG68K_ALU.vhd:266:17  */
  assign n10018_o = n9986_o ? bsout : n10017_o;
  /* TG68K_ALU.vhd:264:17  */
  assign n10019_o = n9985_o ? rot_out : n10018_o;
  /* TG68K_ALU.vhd:261:17  */
  assign n10020_o = n9984_o ? op2out : n10019_o;
  /* TG68K_ALU.vhd:258:17  */
  assign n10021_o = n9982_o ? n9983_o : n10020_o;
  assign n10022_o = n10021_o[7:0];
  /* TG68K_ALU.vhd:256:17  */
  assign n10023_o = n9978_o ? n9981_o : n10022_o;
  assign n10024_o = n10021_o[31:8];
  assign n10025_o = n10166_o[31:8];
  /* TG68K_ALU.vhd:256:17  */
  assign n10026_o = n9978_o ? n10025_o : n10024_o;
  assign n10027_o = {n10026_o, n10023_o};
  /* TG68K_ALU.vhd:254:17  */
  assign n10028_o = n9976_o ? n9977_o : n10027_o;
  /* TG68K_ALU.vhd:252:17  */
  assign n10029_o = n9974_o ? n9975_o : n10028_o;
  /* TG68K_ALU.vhd:241:17  */
  assign n10030_o = n9962_o ? n9973_o : n10029_o;
  /* TG68K_ALU.vhd:226:17  */
  assign n10031_o = n9955_o ? n9959_o : n10030_o;
  assign n10032_o = n10031_o[7:0];
  /* TG68K_ALU.vhd:224:17  */
  assign n10033_o = n9951_o ? n9952_o : n10032_o;
  assign n10034_o = n10031_o[31:8];
  assign n10035_o = n10166_o[31:8];
  /* TG68K_ALU.vhd:224:17  */
  assign n10036_o = n9951_o ? n10035_o : n10034_o;
  /* TG68K_ALU.vhd:293:24  */
  assign n10041_o = exec[29];
  /* TG68K_ALU.vhd:294:34  */
  assign n10042_o = sndopc[11];
  /* TG68K_ALU.vhd:295:51  */
  assign n10043_o = op1out[31];
  /* TG68K_ALU.vhd:295:62  */
  assign n10044_o = op1out[31];
  /* TG68K_ALU.vhd:295:55  */
  assign n10045_o = {n10043_o, n10044_o};
  /* TG68K_ALU.vhd:295:73  */
  assign n10046_o = op1out[31];
  /* TG68K_ALU.vhd:295:66  */
  assign n10047_o = {n10045_o, n10046_o};
  /* TG68K_ALU.vhd:295:84  */
  assign n10048_o = op1out[31:3];
  /* TG68K_ALU.vhd:295:77  */
  assign n10049_o = {n10047_o, n10048_o};
  /* TG68K_ALU.vhd:297:84  */
  assign n10050_o = sndopc[10:9];
  /* TG68K_ALU.vhd:297:77  */
  assign n10052_o = {30'b000000000000000000000000000000, n10050_o};
  /* TG68K_ALU.vhd:294:25  */
  assign n10053_o = n10042_o ? n10049_o : n10052_o;
  /* TG68K_ALU.vhd:293:17  */
  assign n10054_o = n10041_o ? n10053_o : op1out;
  /* TG68K_ALU.vhd:301:24  */
  assign n10055_o = exec[48];
  /* TG68K_ALU.vhd:301:17  */
  assign n10058_o = n10055_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:309:24  */
  assign n10060_o = exec[78];
  /* TG68K_ALU.vhd:310:65  */
  assign n10061_o = op2out[7:4];
  /* TG68K_ALU.vhd:310:57  */
  assign n10063_o = {4'b0000, n10061_o};
  /* TG68K_ALU.vhd:310:78  */
  assign n10065_o = {n10063_o, 4'b0000};
  /* TG68K_ALU.vhd:310:95  */
  assign n10066_o = op2out[3:0];
  /* TG68K_ALU.vhd:310:87  */
  assign n10067_o = {n10065_o, n10066_o};
  /* TG68K_ALU.vhd:311:30  */
  assign n10068_o = ~execopc;
  /* TG68K_ALU.vhd:311:43  */
  assign n10069_o = exec[53];
  /* TG68K_ALU.vhd:311:55  */
  assign n10070_o = ~n10069_o;
  /* TG68K_ALU.vhd:311:35  */
  assign n10071_o = n10070_o & n10068_o;
  /* TG68K_ALU.vhd:311:68  */
  assign n10072_o = exec[29];
  /* TG68K_ALU.vhd:311:82  */
  assign n10073_o = ~n10072_o;
  /* TG68K_ALU.vhd:311:60  */
  assign n10074_o = n10073_o & n10071_o;
  /* TG68K_ALU.vhd:312:38  */
  assign n10075_o = ~long_start;
  /* TG68K_ALU.vhd:312:59  */
  assign n10077_o = exe_datatype == 2'b00;
  /* TG68K_ALU.vhd:312:43  */
  assign n10078_o = n10077_o & n10075_o;
  /* TG68K_ALU.vhd:312:73  */
  assign n10079_o = exec[50];
  /* TG68K_ALU.vhd:312:81  */
  assign n10080_o = ~n10079_o;
  /* TG68K_ALU.vhd:312:65  */
  assign n10081_o = n10080_o & n10078_o;
  /* TG68K_ALU.vhd:314:41  */
  assign n10082_o = ~long_start;
  /* TG68K_ALU.vhd:314:62  */
  assign n10084_o = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:314:46  */
  assign n10085_o = n10084_o & n10082_o;
  /* TG68K_ALU.vhd:314:77  */
  assign n10086_o = exec[47];
  /* TG68K_ALU.vhd:314:93  */
  assign n10087_o = exec[46];
  /* TG68K_ALU.vhd:314:86  */
  assign n10088_o = n10086_o | n10087_o;
  /* TG68K_ALU.vhd:314:103  */
  assign n10089_o = n10088_o | movem_presub;
  /* TG68K_ALU.vhd:314:68  */
  assign n10090_o = n10089_o & n10085_o;
  /* TG68K_ALU.vhd:315:40  */
  assign n10091_o = exec[69];
  /* TG68K_ALU.vhd:315:33  */
  assign n10094_o = n10091_o ? 32'b00000000000000000000000000000110 : 32'b00000000000000000000000000000100;
  /* TG68K_ALU.vhd:314:25  */
  assign n10096_o = n10090_o ? n10094_o : 32'b00000000000000000000000000000010;
  /* TG68K_ALU.vhd:312:25  */
  assign n10098_o = n10081_o ? 32'b00000000000000000000000000000001 : n10096_o;
  /* TG68K_ALU.vhd:324:33  */
  assign n10099_o = exec[28];
  /* TG68K_ALU.vhd:324:59  */
  assign n10100_o = n12945_q[4];
  /* TG68K_ALU.vhd:324:50  */
  assign n10101_o = n10100_o & n10099_o;
  /* TG68K_ALU.vhd:324:75  */
  assign n10102_o = exec[31];
  /* TG68K_ALU.vhd:324:68  */
  assign n10103_o = n10101_o | n10102_o;
  /* TG68K_ALU.vhd:324:25  */
  assign n10105_o = n10103_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:327:41  */
  assign n10106_o = exec[56];
  /* TG68K_ALU.vhd:311:17  */
  assign n10107_o = n10074_o ? n10098_o : op2out;
  /* TG68K_ALU.vhd:311:17  */
  assign n10108_o = n10074_o ? n10058_o : n10106_o;
  /* TG68K_ALU.vhd:311:17  */
  assign n10109_o = n10074_o ? 1'b0 : n10105_o;
  assign n10110_o = n10107_o[15:0];
  /* TG68K_ALU.vhd:309:17  */
  assign n10111_o = n10060_o ? n10067_o : n10110_o;
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n10112_o = n10107_o[31:16];
  /* TG68KdotC_Kernel.vhd:1401:33  */
  assign n10113_o = op2out[31:16];
  /* TG68K_ALU.vhd:309:17  */
  assign n10114_o = n10060_o ? n10113_o : n10112_o;
  /* TG68K_ALU.vhd:309:17  */
  assign n10116_o = n10060_o ? n10058_o : n10108_o;
  /* TG68K_ALU.vhd:309:17  */
  assign n10117_o = n10060_o ? 1'b0 : n10109_o;
  /* TG68K_ALU.vhd:331:24  */
  assign n10118_o = exec[69];
  /* TG68K_ALU.vhd:331:43  */
  assign n10119_o = n10118_o | check_aligned;
  /* TG68K_ALU.vhd:332:36  */
  assign n10120_o = ~movem_presub;
  /* TG68K_ALU.vhd:333:64  */
  assign n10121_o = ~long_start;
  /* TG68K_ALU.vhd:333:48  */
  assign n10122_o = n10121_o & non_aligned;
  /* TG68KdotC_Kernel.vhd:1275:33  */
  assign n10124_o = {n10114_o, n10111_o};
  /* TG68K_ALU.vhd:333:25  */
  assign n10125_o = n10122_o ? 32'b00000000000000000000000000000000 : n10124_o;
  /* TG68K_ALU.vhd:337:64  */
  assign n10126_o = ~long_start;
  /* TG68K_ALU.vhd:337:48  */
  assign n10127_o = n10126_o & non_aligned;
  /* TG68K_ALU.vhd:338:44  */
  assign n10129_o = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:338:27  */
  assign n10132_o = n10129_o ? 32'b00000000000000000000000000001000 : 32'b00000000000000000000000000000100;
  assign n10133_o = {n10114_o, n10111_o};
  /* TG68K_ALU.vhd:337:25  */
  assign n10134_o = n10127_o ? n10132_o : n10133_o;
  /* TG68K_ALU.vhd:332:19  */
  assign n10135_o = n10120_o ? n10125_o : n10134_o;
  assign n10136_o = {n10114_o, n10111_o};
  /* TG68K_ALU.vhd:331:17  */
  assign n10137_o = n10119_o ? n10135_o : n10136_o;
  /* TG68K_ALU.vhd:347:28  */
  assign n10138_o = ~opaddsub;
  /* TG68K_ALU.vhd:347:33  */
  assign n10139_o = n10138_o | long_start;
  /* TG68K_ALU.vhd:348:43  */
  assign n10141_o = {1'b0, addsub_b};
  /* TG68K_ALU.vhd:348:57  */
  assign n10142_o = c_in[0];
  /* TG68K_ALU.vhd:348:52  */
  assign n10143_o = {n10141_o, n10142_o};
  /* TG68K_ALU.vhd:350:48  */
  assign n10145_o = {1'b0, addsub_b};
  /* TG68K_ALU.vhd:350:62  */
  assign n10146_o = c_in[0];
  /* TG68K_ALU.vhd:350:57  */
  assign n10147_o = {n10145_o, n10146_o};
  /* TG68K_ALU.vhd:350:40  */
  assign n10148_o = ~n10147_o;
  /* TG68K_ALU.vhd:347:17  */
  assign n10149_o = n10139_o ? n10143_o : n10148_o;
  /* TG68K_ALU.vhd:352:36  */
  assign n10151_o = {1'b0, addsub_a};
  /* TG68K_ALU.vhd:352:57  */
  assign n10152_o = notaddsub_b[0];
  /* TG68K_ALU.vhd:352:45  */
  assign n10153_o = {n10151_o, n10152_o};
  /* TG68K_ALU.vhd:352:61  */
  assign n10154_o = n10153_o + notaddsub_b;
  /* TG68K_ALU.vhd:353:38  */
  assign n10155_o = add_result[9];
  /* TG68K_ALU.vhd:353:54  */
  assign n10156_o = addsub_a[8];
  /* TG68K_ALU.vhd:353:42  */
  assign n10157_o = n10155_o ^ n10156_o;
  /* TG68K_ALU.vhd:353:70  */
  assign n10158_o = addsub_b[8];
  /* TG68K_ALU.vhd:353:58  */
  assign n10159_o = n10157_o ^ n10158_o;
  /* TG68K_ALU.vhd:354:38  */
  assign n10160_o = add_result[17];
  /* TG68K_ALU.vhd:354:55  */
  assign n10161_o = addsub_a[16];
  /* TG68K_ALU.vhd:354:43  */
  assign n10162_o = n10160_o ^ n10161_o;
  /* TG68K_ALU.vhd:354:72  */
  assign n10163_o = addsub_b[16];
  /* TG68K_ALU.vhd:354:60  */
  assign n10164_o = n10162_o ^ n10163_o;
  /* TG68K_ALU.vhd:355:38  */
  assign n10165_o = add_result[33];
  /* TG68K_ALU.vhd:356:39  */
  assign n10166_o = add_result[32:1];
  /* TG68K_ALU.vhd:357:39  */
  assign n10167_o = c_in[1];
  /* TG68K_ALU.vhd:357:57  */
  assign n10168_o = add_result[8];
  /* TG68K_ALU.vhd:357:43  */
  assign n10169_o = n10167_o ^ n10168_o;
  /* TG68K_ALU.vhd:357:73  */
  assign n10170_o = addsub_a[7];
  /* TG68K_ALU.vhd:357:61  */
  assign n10171_o = n10169_o ^ n10170_o;
  /* TG68K_ALU.vhd:357:89  */
  assign n10172_o = addsub_b[7];
  /* TG68K_ALU.vhd:357:77  */
  assign n10173_o = n10171_o ^ n10172_o;
  /* TG68K_ALU.vhd:358:39  */
  assign n10174_o = c_in[2];
  /* TG68K_ALU.vhd:358:57  */
  assign n10175_o = add_result[16];
  /* TG68K_ALU.vhd:358:43  */
  assign n10176_o = n10174_o ^ n10175_o;
  /* TG68K_ALU.vhd:358:74  */
  assign n10177_o = addsub_a[15];
  /* TG68K_ALU.vhd:358:62  */
  assign n10178_o = n10176_o ^ n10177_o;
  /* TG68K_ALU.vhd:358:91  */
  assign n10179_o = addsub_b[15];
  /* TG68K_ALU.vhd:358:79  */
  assign n10180_o = n10178_o ^ n10179_o;
  /* TG68K_ALU.vhd:359:39  */
  assign n10181_o = c_in[3];
  /* TG68K_ALU.vhd:359:57  */
  assign n10182_o = add_result[32];
  /* TG68K_ALU.vhd:359:43  */
  assign n10183_o = n10181_o ^ n10182_o;
  /* TG68K_ALU.vhd:359:74  */
  assign n10184_o = addsub_a[31];
  /* TG68K_ALU.vhd:359:62  */
  assign n10185_o = n10183_o ^ n10184_o;
  /* TG68K_ALU.vhd:359:91  */
  assign n10186_o = addsub_b[31];
  /* TG68K_ALU.vhd:359:79  */
  assign n10187_o = n10185_o ^ n10186_o;
  /* TG68K_ALU.vhd:360:30  */
  assign n10188_o = c_in[3:1];
  /* TG68K_ALU.vhd:370:32  */
  assign n10192_o = c_in[1];
  /* TG68K_ALU.vhd:370:46  */
  assign n10193_o = add_result[8:0];
  /* TG68K_ALU.vhd:370:35  */
  assign n10194_o = {n10192_o, n10193_o};
  /* TG68K_ALU.vhd:372:38  */
  assign n10195_o = op1out[4];
  /* TG68K_ALU.vhd:372:52  */
  assign n10196_o = op2out[4];
  /* TG68K_ALU.vhd:372:42  */
  assign n10197_o = n10195_o ^ n10196_o;
  /* TG68K_ALU.vhd:372:67  */
  assign n10198_o = bcd_pur[5];
  /* TG68K_ALU.vhd:372:56  */
  assign n10199_o = n10197_o ^ n10198_o;
  /* TG68K_ALU.vhd:373:17  */
  assign n10202_o = halve_carry ? 4'b0110 : 4'b0000;
  /* TG68K_ALU.vhd:376:27  */
  assign n10205_o = bcd_pur[9];
  assign n10207_o = n10203_o[7:4];
  /* TG68K_ALU.vhd:376:17  */
  assign n10208_o = n10205_o ? 4'b0110 : n10207_o;
  assign n10209_o = n10203_o[8];
  /* TG68K_ALU.vhd:379:24  */
  assign n10210_o = exec[12];
  /* TG68K_ALU.vhd:380:47  */
  assign n10211_o = bcd_pur[8];
  /* TG68K_ALU.vhd:380:36  */
  assign n10212_o = ~n10211_o;
  /* TG68K_ALU.vhd:380:60  */
  assign n10213_o = bcd_a[7];
  /* TG68K_ALU.vhd:380:51  */
  assign n10214_o = n10212_o & n10213_o;
  /* TG68K_ALU.vhd:382:41  */
  assign n10215_o = bcd_pur[9:1];
  /* TG68K_ALU.vhd:382:54  */
  assign n10216_o = n10215_o + bcd_kor;
  /* TG68K_ALU.vhd:383:36  */
  assign n10217_o = bcd_pur[4];
  /* TG68K_ALU.vhd:383:52  */
  assign n10218_o = bcd_pur[3];
  /* TG68K_ALU.vhd:383:66  */
  assign n10219_o = bcd_pur[2];
  /* TG68K_ALU.vhd:383:56  */
  assign n10220_o = n10218_o | n10219_o;
  /* TG68K_ALU.vhd:383:40  */
  assign n10221_o = n10217_o & n10220_o;
  /* TG68K_ALU.vhd:383:25  */
  assign n10223_o = n10221_o ? 4'b0110 : n10202_o;
  /* TG68K_ALU.vhd:386:36  */
  assign n10224_o = bcd_pur[8];
  /* TG68K_ALU.vhd:386:52  */
  assign n10225_o = bcd_pur[7];
  /* TG68K_ALU.vhd:386:66  */
  assign n10226_o = bcd_pur[6];
  /* TG68K_ALU.vhd:386:56  */
  assign n10227_o = n10225_o | n10226_o;
  /* TG68K_ALU.vhd:386:81  */
  assign n10228_o = bcd_pur[5];
  /* TG68K_ALU.vhd:386:96  */
  assign n10229_o = bcd_pur[4];
  /* TG68K_ALU.vhd:386:85  */
  assign n10230_o = n10228_o & n10229_o;
  /* TG68K_ALU.vhd:386:112  */
  assign n10231_o = bcd_pur[3];
  /* TG68K_ALU.vhd:386:126  */
  assign n10232_o = bcd_pur[2];
  /* TG68K_ALU.vhd:386:116  */
  assign n10233_o = n10231_o | n10232_o;
  /* TG68K_ALU.vhd:386:100  */
  assign n10234_o = n10230_o & n10233_o;
  /* TG68K_ALU.vhd:386:70  */
  assign n10235_o = n10227_o | n10234_o;
  /* TG68K_ALU.vhd:386:40  */
  assign n10236_o = n10224_o & n10235_o;
  /* TG68K_ALU.vhd:386:25  */
  assign n10238_o = n10236_o ? 4'b0110 : n10208_o;
  /* TG68K_ALU.vhd:390:43  */
  assign n10239_o = bcd_pur[8];
  /* TG68K_ALU.vhd:390:60  */
  assign n10240_o = bcd_a[7];
  /* TG68K_ALU.vhd:390:51  */
  assign n10241_o = ~n10240_o;
  /* TG68K_ALU.vhd:390:47  */
  assign n10242_o = n10239_o & n10241_o;
  /* TG68K_ALU.vhd:392:41  */
  assign n10243_o = bcd_pur[9:1];
  /* TG68K_ALU.vhd:392:54  */
  assign n10244_o = n10243_o - bcd_kor;
  assign n10245_o = {n10238_o, n10223_o};
  assign n10246_o = {n10208_o, n10202_o};
  /* TG68K_ALU.vhd:379:17  */
  assign n10247_o = n10210_o ? n10245_o : n10246_o;
  /* TG68K_ALU.vhd:379:17  */
  assign n10248_o = n10210_o ? n10214_o : n10242_o;
  /* TG68K_ALU.vhd:379:17  */
  assign n10249_o = n10210_o ? n10216_o : n10244_o;
  /* TG68K_ALU.vhd:394:23  */
  assign n10250_o = cpu[1];
  /* TG68K_ALU.vhd:394:17  */
  assign n10252_o = n10250_o ? 1'b0 : n10248_o;
  /* TG68K_ALU.vhd:397:39  */
  assign n10253_o = bcd_pur[9];
  /* TG68K_ALU.vhd:397:51  */
  assign n10254_o = bcd_a[8];
  /* TG68K_ALU.vhd:397:43  */
  assign n10255_o = n10253_o | n10254_o;
  /* TG68K_ALU.vhd:409:44  */
  assign n10260_o = opcode[7:6];
  /* TG68K_ALU.vhd:410:41  */
  assign n10262_o = n10260_o == 2'b01;
  /* TG68K_ALU.vhd:412:41  */
  assign n10264_o = n10260_o == 2'b11;
  assign n10265_o = {n10264_o, n10262_o};
  /* TG68K_ALU.vhd:409:33  */
  always @*
    case (n10265_o)
      2'b10: n10268_o = 1'b0;
      2'b01: n10268_o = 1'b1;
      default: n10268_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:409:33  */
  always @*
    case (n10265_o)
      2'b10: n10272_o = 1'b1;
      2'b01: n10272_o = 1'b0;
      default: n10272_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:419:30  */
  assign n10278_o = exe_opcode[8];
  /* TG68K_ALU.vhd:419:33  */
  assign n10279_o = ~n10278_o;
  /* TG68K_ALU.vhd:420:38  */
  assign n10280_o = exe_opcode[5:4];
  /* TG68K_ALU.vhd:420:50  */
  assign n10282_o = n10280_o == 2'b00;
  /* TG68K_ALU.vhd:421:53  */
  assign n10283_o = sndopc[4:0];
  /* TG68K_ALU.vhd:423:58  */
  assign n10284_o = sndopc[2:0];
  /* TG68K_ALU.vhd:423:51  */
  assign n10286_o = {2'b00, n10284_o};
  /* TG68K_ALU.vhd:420:25  */
  assign n10287_o = n10282_o ? n10283_o : n10286_o;
  /* TG68K_ALU.vhd:426:38  */
  assign n10288_o = exe_opcode[5:4];
  /* TG68K_ALU.vhd:426:50  */
  assign n10290_o = n10288_o == 2'b00;
  /* TG68K_ALU.vhd:427:53  */
  assign n10291_o = reg_qb[4:0];
  /* TG68K_ALU.vhd:429:58  */
  assign n10292_o = reg_qb[2:0];
  /* TG68K_ALU.vhd:429:51  */
  assign n10294_o = {2'b00, n10292_o};
  /* TG68K_ALU.vhd:426:25  */
  assign n10295_o = n10290_o ? n10291_o : n10294_o;
  /* TG68K_ALU.vhd:419:17  */
  assign n10296_o = n10279_o ? n10287_o : n10295_o;
  /* TG68K_ALU.vhd:435:65  */
  assign n10302_o = ~one_bit_in;
  /* TG68K_ALU.vhd:435:61  */
  assign n10303_o = bchg & n10302_o;
  /* TG68K_ALU.vhd:435:81  */
  assign n10304_o = n10303_o | bset;
  /* TG68K_ALU.vhd:456:42  */
  assign n10310_o = opcode[5:4];
  /* TG68K_ALU.vhd:456:55  */
  assign n10312_o = n10310_o == 2'b00;
  /* TG68K_ALU.vhd:456:33  */
  assign n10315_o = n10312_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:459:44  */
  assign n10317_o = opcode[10:8];
  /* TG68K_ALU.vhd:460:41  */
  assign n10319_o = n10317_o == 3'b010;
  /* TG68K_ALU.vhd:461:41  */
  assign n10321_o = n10317_o == 3'b011;
  /* TG68K_ALU.vhd:463:41  */
  assign n10323_o = n10317_o == 3'b101;
  /* TG68K_ALU.vhd:464:41  */
  assign n10325_o = n10317_o == 3'b110;
  /* TG68K_ALU.vhd:465:41  */
  assign n10327_o = n10317_o == 3'b111;
  assign n10328_o = {n10327_o, n10325_o, n10323_o, n10321_o, n10319_o};
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10328_o)
      5'b10000: n10331_o = 1'b0;
      5'b01000: n10331_o = 1'b1;
      5'b00100: n10331_o = 1'b0;
      5'b00010: n10331_o = 1'b0;
      5'b00001: n10331_o = 1'b0;
      default: n10331_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10328_o)
      5'b10000: n10335_o = 1'b0;
      5'b01000: n10335_o = 1'b0;
      5'b00100: n10335_o = 1'b0;
      5'b00010: n10335_o = 1'b0;
      5'b00001: n10335_o = 1'b1;
      default: n10335_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10328_o)
      5'b10000: n10339_o = 1'b1;
      5'b01000: n10339_o = 1'b0;
      5'b00100: n10339_o = 1'b0;
      5'b00010: n10339_o = 1'b0;
      5'b00001: n10339_o = 1'b0;
      default: n10339_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10328_o)
      5'b10000: n10343_o = 1'b0;
      5'b01000: n10343_o = 1'b0;
      5'b00100: n10343_o = 1'b0;
      5'b00010: n10343_o = 1'b1;
      5'b00001: n10343_o = 1'b0;
      default: n10343_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10328_o)
      5'b10000: n10347_o = 1'b0;
      5'b01000: n10347_o = 1'b0;
      5'b00100: n10347_o = 1'b1;
      5'b00010: n10347_o = 1'b0;
      5'b00001: n10347_o = 1'b0;
      default: n10347_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10328_o)
      5'b10000: n10350_o = 1'b1;
      5'b01000: n10350_o = n10315_o;
      5'b00100: n10350_o = n10315_o;
      5'b00010: n10350_o = n10315_o;
      5'b00001: n10350_o = n10315_o;
      default: n10350_o = n10315_o;
    endcase
  /* TG68K_ALU.vhd:469:42  */
  assign n10351_o = opcode[4:3];
  /* TG68K_ALU.vhd:469:54  */
  assign n10353_o = n10351_o == 2'b00;
  /* TG68K_ALU.vhd:469:33  */
  assign n10356_o = n10353_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:472:53  */
  assign n10358_o = result[39:32];
  /* TG68K_ALU.vhd:490:38  */
  assign n10376_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10378_o = $unsigned(5'b00000) > $unsigned(n10376_o);
  assign n10381_o = reg_qb[0];
  assign n10382_o = bf_set2[0];
  /* TG68K_ALU.vhd:476:17  */
  assign n10383_o = bf_ins ? n10381_o : n10382_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10384_o = n10378_o ? 1'b0 : n10383_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10389_o = n10378_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:490:38  */
  assign n10392_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10394_o = $unsigned(5'b00001) > $unsigned(n10392_o);
  assign n10397_o = reg_qb[1];
  assign n10398_o = bf_set2[1];
  /* TG68K_ALU.vhd:476:17  */
  assign n10399_o = bf_ins ? n10397_o : n10398_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10400_o = n10394_o ? 1'b0 : n10399_o;
  assign n10404_o = n10390_o[1];
  /* TG68K_ALU.vhd:490:25  */
  assign n10405_o = n10394_o ? 1'b1 : n10404_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10407_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10409_o = $unsigned(5'b00010) > $unsigned(n10407_o);
  assign n10412_o = reg_qb[2];
  assign n10413_o = bf_set2[2];
  /* TG68K_ALU.vhd:476:17  */
  assign n10414_o = bf_ins ? n10412_o : n10413_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10415_o = n10409_o ? 1'b0 : n10414_o;
  assign n10419_o = n10390_o[2];
  /* TG68K_ALU.vhd:490:25  */
  assign n10420_o = n10409_o ? 1'b1 : n10419_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10422_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10424_o = $unsigned(5'b00011) > $unsigned(n10422_o);
  assign n10427_o = reg_qb[3];
  assign n10428_o = bf_set2[3];
  /* TG68K_ALU.vhd:476:17  */
  assign n10429_o = bf_ins ? n10427_o : n10428_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10430_o = n10424_o ? 1'b0 : n10429_o;
  assign n10434_o = n10390_o[3];
  /* TG68K_ALU.vhd:490:25  */
  assign n10435_o = n10424_o ? 1'b1 : n10434_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10437_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10439_o = $unsigned(5'b00100) > $unsigned(n10437_o);
  assign n10442_o = reg_qb[4];
  assign n10443_o = bf_set2[4];
  /* TG68K_ALU.vhd:476:17  */
  assign n10444_o = bf_ins ? n10442_o : n10443_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10445_o = n10439_o ? 1'b0 : n10444_o;
  assign n10449_o = n10390_o[4];
  /* TG68K_ALU.vhd:490:25  */
  assign n10450_o = n10439_o ? 1'b1 : n10449_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10452_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10454_o = $unsigned(5'b00101) > $unsigned(n10452_o);
  assign n10457_o = reg_qb[5];
  assign n10458_o = bf_set2[5];
  /* TG68K_ALU.vhd:476:17  */
  assign n10459_o = bf_ins ? n10457_o : n10458_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10460_o = n10454_o ? 1'b0 : n10459_o;
  assign n10464_o = n10390_o[5];
  /* TG68K_ALU.vhd:490:25  */
  assign n10465_o = n10454_o ? 1'b1 : n10464_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10467_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10469_o = $unsigned(5'b00110) > $unsigned(n10467_o);
  assign n10472_o = reg_qb[6];
  assign n10473_o = bf_set2[6];
  /* TG68K_ALU.vhd:476:17  */
  assign n10474_o = bf_ins ? n10472_o : n10473_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10475_o = n10469_o ? 1'b0 : n10474_o;
  assign n10479_o = n10390_o[6];
  /* TG68K_ALU.vhd:490:25  */
  assign n10480_o = n10469_o ? 1'b1 : n10479_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10482_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10484_o = $unsigned(5'b00111) > $unsigned(n10482_o);
  assign n10487_o = reg_qb[7];
  assign n10488_o = bf_set2[7];
  /* TG68K_ALU.vhd:476:17  */
  assign n10489_o = bf_ins ? n10487_o : n10488_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10490_o = n10484_o ? 1'b0 : n10489_o;
  assign n10494_o = n10390_o[7];
  /* TG68K_ALU.vhd:490:25  */
  assign n10495_o = n10484_o ? 1'b1 : n10494_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10497_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10499_o = $unsigned(5'b01000) > $unsigned(n10497_o);
  assign n10502_o = reg_qb[8];
  assign n10503_o = bf_set2[8];
  /* TG68K_ALU.vhd:476:17  */
  assign n10504_o = bf_ins ? n10502_o : n10503_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10505_o = n10499_o ? 1'b0 : n10504_o;
  assign n10509_o = n10390_o[8];
  /* TG68K_ALU.vhd:490:25  */
  assign n10510_o = n10499_o ? 1'b1 : n10509_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10512_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10514_o = $unsigned(5'b01001) > $unsigned(n10512_o);
  assign n10517_o = reg_qb[9];
  assign n10518_o = bf_set2[9];
  /* TG68K_ALU.vhd:476:17  */
  assign n10519_o = bf_ins ? n10517_o : n10518_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10520_o = n10514_o ? 1'b0 : n10519_o;
  assign n10524_o = n10390_o[9];
  /* TG68K_ALU.vhd:490:25  */
  assign n10525_o = n10514_o ? 1'b1 : n10524_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10527_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10529_o = $unsigned(5'b01010) > $unsigned(n10527_o);
  assign n10532_o = reg_qb[10];
  assign n10533_o = bf_set2[10];
  /* TG68K_ALU.vhd:476:17  */
  assign n10534_o = bf_ins ? n10532_o : n10533_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10535_o = n10529_o ? 1'b0 : n10534_o;
  assign n10539_o = n10390_o[10];
  /* TG68K_ALU.vhd:490:25  */
  assign n10540_o = n10529_o ? 1'b1 : n10539_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10542_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10544_o = $unsigned(5'b01011) > $unsigned(n10542_o);
  assign n10547_o = reg_qb[11];
  assign n10548_o = bf_set2[11];
  /* TG68K_ALU.vhd:476:17  */
  assign n10549_o = bf_ins ? n10547_o : n10548_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10550_o = n10544_o ? 1'b0 : n10549_o;
  assign n10554_o = n10390_o[11];
  /* TG68K_ALU.vhd:490:25  */
  assign n10555_o = n10544_o ? 1'b1 : n10554_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10557_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10559_o = $unsigned(5'b01100) > $unsigned(n10557_o);
  assign n10562_o = reg_qb[12];
  assign n10563_o = bf_set2[12];
  /* TG68K_ALU.vhd:476:17  */
  assign n10564_o = bf_ins ? n10562_o : n10563_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10565_o = n10559_o ? 1'b0 : n10564_o;
  assign n10569_o = n10390_o[12];
  /* TG68K_ALU.vhd:490:25  */
  assign n10570_o = n10559_o ? 1'b1 : n10569_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10572_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10574_o = $unsigned(5'b01101) > $unsigned(n10572_o);
  assign n10577_o = reg_qb[13];
  assign n10578_o = bf_set2[13];
  /* TG68K_ALU.vhd:476:17  */
  assign n10579_o = bf_ins ? n10577_o : n10578_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10580_o = n10574_o ? 1'b0 : n10579_o;
  assign n10584_o = n10390_o[13];
  /* TG68K_ALU.vhd:490:25  */
  assign n10585_o = n10574_o ? 1'b1 : n10584_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10587_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10589_o = $unsigned(5'b01110) > $unsigned(n10587_o);
  assign n10592_o = reg_qb[14];
  assign n10593_o = bf_set2[14];
  /* TG68K_ALU.vhd:476:17  */
  assign n10594_o = bf_ins ? n10592_o : n10593_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10595_o = n10589_o ? 1'b0 : n10594_o;
  assign n10599_o = n10390_o[14];
  /* TG68K_ALU.vhd:490:25  */
  assign n10600_o = n10589_o ? 1'b1 : n10599_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10602_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10604_o = $unsigned(5'b01111) > $unsigned(n10602_o);
  assign n10607_o = reg_qb[15];
  assign n10608_o = bf_set2[15];
  /* TG68K_ALU.vhd:476:17  */
  assign n10609_o = bf_ins ? n10607_o : n10608_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10610_o = n10604_o ? 1'b0 : n10609_o;
  assign n10614_o = n10390_o[15];
  /* TG68K_ALU.vhd:490:25  */
  assign n10615_o = n10604_o ? 1'b1 : n10614_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10617_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10619_o = $unsigned(5'b10000) > $unsigned(n10617_o);
  assign n10622_o = reg_qb[16];
  assign n10623_o = bf_set2[16];
  /* TG68K_ALU.vhd:476:17  */
  assign n10624_o = bf_ins ? n10622_o : n10623_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10625_o = n10619_o ? 1'b0 : n10624_o;
  assign n10629_o = n10390_o[16];
  /* TG68K_ALU.vhd:490:25  */
  assign n10630_o = n10619_o ? 1'b1 : n10629_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10632_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10634_o = $unsigned(5'b10001) > $unsigned(n10632_o);
  assign n10637_o = reg_qb[17];
  assign n10638_o = bf_set2[17];
  /* TG68K_ALU.vhd:476:17  */
  assign n10639_o = bf_ins ? n10637_o : n10638_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10640_o = n10634_o ? 1'b0 : n10639_o;
  assign n10644_o = n10390_o[17];
  /* TG68K_ALU.vhd:490:25  */
  assign n10645_o = n10634_o ? 1'b1 : n10644_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10647_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10649_o = $unsigned(5'b10010) > $unsigned(n10647_o);
  assign n10652_o = reg_qb[18];
  assign n10653_o = bf_set2[18];
  /* TG68K_ALU.vhd:476:17  */
  assign n10654_o = bf_ins ? n10652_o : n10653_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10655_o = n10649_o ? 1'b0 : n10654_o;
  assign n10659_o = n10390_o[18];
  /* TG68K_ALU.vhd:490:25  */
  assign n10660_o = n10649_o ? 1'b1 : n10659_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10662_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10664_o = $unsigned(5'b10011) > $unsigned(n10662_o);
  assign n10667_o = reg_qb[19];
  assign n10668_o = bf_set2[19];
  /* TG68K_ALU.vhd:476:17  */
  assign n10669_o = bf_ins ? n10667_o : n10668_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10670_o = n10664_o ? 1'b0 : n10669_o;
  assign n10674_o = n10390_o[19];
  /* TG68K_ALU.vhd:490:25  */
  assign n10675_o = n10664_o ? 1'b1 : n10674_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10677_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10679_o = $unsigned(5'b10100) > $unsigned(n10677_o);
  assign n10682_o = reg_qb[20];
  assign n10683_o = bf_set2[20];
  /* TG68K_ALU.vhd:476:17  */
  assign n10684_o = bf_ins ? n10682_o : n10683_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10685_o = n10679_o ? 1'b0 : n10684_o;
  assign n10689_o = n10390_o[20];
  /* TG68K_ALU.vhd:490:25  */
  assign n10690_o = n10679_o ? 1'b1 : n10689_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10692_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10694_o = $unsigned(5'b10101) > $unsigned(n10692_o);
  assign n10697_o = reg_qb[21];
  assign n10698_o = bf_set2[21];
  /* TG68K_ALU.vhd:476:17  */
  assign n10699_o = bf_ins ? n10697_o : n10698_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10700_o = n10694_o ? 1'b0 : n10699_o;
  assign n10704_o = n10390_o[21];
  /* TG68K_ALU.vhd:490:25  */
  assign n10705_o = n10694_o ? 1'b1 : n10704_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10707_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10709_o = $unsigned(5'b10110) > $unsigned(n10707_o);
  assign n10712_o = reg_qb[22];
  assign n10713_o = bf_set2[22];
  /* TG68K_ALU.vhd:476:17  */
  assign n10714_o = bf_ins ? n10712_o : n10713_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10715_o = n10709_o ? 1'b0 : n10714_o;
  assign n10719_o = n10390_o[22];
  /* TG68K_ALU.vhd:490:25  */
  assign n10720_o = n10709_o ? 1'b1 : n10719_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10722_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10724_o = $unsigned(5'b10111) > $unsigned(n10722_o);
  assign n10727_o = reg_qb[23];
  assign n10728_o = bf_set2[23];
  /* TG68K_ALU.vhd:476:17  */
  assign n10729_o = bf_ins ? n10727_o : n10728_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10730_o = n10724_o ? 1'b0 : n10729_o;
  assign n10734_o = n10390_o[23];
  /* TG68K_ALU.vhd:490:25  */
  assign n10735_o = n10724_o ? 1'b1 : n10734_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10737_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10739_o = $unsigned(5'b11000) > $unsigned(n10737_o);
  assign n10742_o = reg_qb[24];
  assign n10743_o = bf_set2[24];
  /* TG68K_ALU.vhd:476:17  */
  assign n10744_o = bf_ins ? n10742_o : n10743_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10745_o = n10739_o ? 1'b0 : n10744_o;
  assign n10749_o = n10390_o[24];
  /* TG68K_ALU.vhd:490:25  */
  assign n10750_o = n10739_o ? 1'b1 : n10749_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10752_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10754_o = $unsigned(5'b11001) > $unsigned(n10752_o);
  assign n10757_o = reg_qb[25];
  assign n10758_o = bf_set2[25];
  /* TG68K_ALU.vhd:476:17  */
  assign n10759_o = bf_ins ? n10757_o : n10758_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10760_o = n10754_o ? 1'b0 : n10759_o;
  assign n10764_o = n10390_o[25];
  /* TG68K_ALU.vhd:490:25  */
  assign n10765_o = n10754_o ? 1'b1 : n10764_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10767_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10769_o = $unsigned(5'b11010) > $unsigned(n10767_o);
  assign n10772_o = reg_qb[26];
  assign n10773_o = bf_set2[26];
  /* TG68K_ALU.vhd:476:17  */
  assign n10774_o = bf_ins ? n10772_o : n10773_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10775_o = n10769_o ? 1'b0 : n10774_o;
  assign n10779_o = n10390_o[26];
  /* TG68K_ALU.vhd:490:25  */
  assign n10780_o = n10769_o ? 1'b1 : n10779_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10782_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10784_o = $unsigned(5'b11011) > $unsigned(n10782_o);
  assign n10787_o = reg_qb[27];
  assign n10788_o = bf_set2[27];
  /* TG68K_ALU.vhd:476:17  */
  assign n10789_o = bf_ins ? n10787_o : n10788_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10790_o = n10784_o ? 1'b0 : n10789_o;
  assign n10794_o = n10390_o[27];
  /* TG68K_ALU.vhd:490:25  */
  assign n10795_o = n10784_o ? 1'b1 : n10794_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10797_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10799_o = $unsigned(5'b11100) > $unsigned(n10797_o);
  assign n10802_o = reg_qb[28];
  assign n10803_o = bf_set2[28];
  /* TG68K_ALU.vhd:476:17  */
  assign n10804_o = bf_ins ? n10802_o : n10803_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10805_o = n10799_o ? 1'b0 : n10804_o;
  assign n10809_o = n10390_o[28];
  /* TG68K_ALU.vhd:490:25  */
  assign n10810_o = n10799_o ? 1'b1 : n10809_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10812_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10814_o = $unsigned(5'b11101) > $unsigned(n10812_o);
  assign n10817_o = reg_qb[29];
  assign n10818_o = bf_set2[29];
  /* TG68K_ALU.vhd:476:17  */
  assign n10819_o = bf_ins ? n10817_o : n10818_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10820_o = n10814_o ? 1'b0 : n10819_o;
  assign n10824_o = n10390_o[29];
  /* TG68K_ALU.vhd:490:25  */
  assign n10825_o = n10814_o ? 1'b1 : n10824_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10827_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10829_o = $unsigned(5'b11110) > $unsigned(n10827_o);
  assign n10832_o = reg_qb[30];
  assign n10833_o = bf_set2[30];
  /* TG68K_ALU.vhd:476:17  */
  assign n10834_o = bf_ins ? n10832_o : n10833_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10835_o = n10829_o ? 1'b0 : n10834_o;
  assign n10836_o = reg_qb[31];
  assign n10837_o = bf_set2[31];
  /* TG68K_ALU.vhd:476:17  */
  assign n10838_o = bf_ins ? n10836_o : n10837_o;
  assign n10839_o = n10390_o[30];
  /* TG68K_ALU.vhd:490:25  */
  assign n10840_o = n10829_o ? 1'b1 : n10839_o;
  assign n10841_o = n10390_o[31];
  /* TG68K_ALU.vhd:490:38  */
  assign n10842_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10844_o = $unsigned(5'b11111) > $unsigned(n10842_o);
  /* TG68K_ALU.vhd:490:25  */
  assign n10847_o = n10844_o ? 1'b0 : n10838_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10848_o = n10844_o ? 1'b1 : n10841_o;
  /* TG68K_ALU.vhd:496:37  */
  assign n10850_o = bf_width[4:0];  // trunc
  /* TG68K_ALU.vhd:497:32  */
  assign n10853_o = bf_nflag & bf_exts;
  /* TG68K_ALU.vhd:498:47  */
  assign n10854_o = datareg | unshifted_bitmask;
  /* TG68K_ALU.vhd:497:17  */
  assign n10855_o = n10853_o ? n10854_o : datareg;
  /* TG68K_ALU.vhd:504:30  */
  assign n10856_o = bf_loffset[4];
  /* TG68K_ALU.vhd:505:57  */
  assign n10857_o = unshifted_bitmask[15:0];
  /* TG68K_ALU.vhd:505:88  */
  assign n10858_o = unshifted_bitmask[31:16];
  /* TG68K_ALU.vhd:505:70  */
  assign n10859_o = {n10857_o, n10858_o};
  /* TG68K_ALU.vhd:504:17  */
  assign n10860_o = n10856_o ? n10859_o : unshifted_bitmask;
  /* TG68K_ALU.vhd:509:30  */
  assign n10861_o = bf_loffset[3];
  /* TG68K_ALU.vhd:510:64  */
  assign n10862_o = bitmaskmux3[23:0];
  /* TG68K_ALU.vhd:510:89  */
  assign n10863_o = bitmaskmux3[31:24];
  /* TG68K_ALU.vhd:510:77  */
  assign n10864_o = {n10862_o, n10863_o};
  /* TG68K_ALU.vhd:509:17  */
  assign n10865_o = n10861_o ? n10864_o : bitmaskmux3;
  /* TG68K_ALU.vhd:514:30  */
  assign n10866_o = bf_loffset[2];
  /* TG68K_ALU.vhd:515:51  */
  assign n10868_o = {bitmaskmux2, 4'b1111};
  /* TG68K_ALU.vhd:517:71  */
  assign n10869_o = bitmaskmux2[31:28];
  assign n10870_o = n10868_o[3:0];
  /* TG68K_ALU.vhd:516:25  */
  assign n10871_o = bf_d32 ? n10869_o : n10870_o;
  assign n10872_o = n10868_o[35:4];
  /* TG68K_ALU.vhd:520:46  */
  assign n10874_o = {4'b1111, bitmaskmux2};
  assign n10875_o = {n10872_o, n10871_o};
  /* TG68K_ALU.vhd:514:17  */
  assign n10876_o = n10866_o ? n10875_o : n10874_o;
  /* TG68K_ALU.vhd:522:30  */
  assign n10877_o = bf_loffset[1];
  /* TG68K_ALU.vhd:523:51  */
  assign n10879_o = {bitmaskmux1, 2'b11};
  /* TG68K_ALU.vhd:525:71  */
  assign n10880_o = bitmaskmux1[31:30];
  assign n10881_o = n10879_o[1:0];
  /* TG68K_ALU.vhd:524:25  */
  assign n10882_o = bf_d32 ? n10880_o : n10881_o;
  assign n10883_o = n10879_o[37:2];
  /* TG68K_ALU.vhd:528:44  */
  assign n10885_o = {2'b11, bitmaskmux1};
  assign n10886_o = {n10883_o, n10882_o};
  /* TG68K_ALU.vhd:522:17  */
  assign n10887_o = n10877_o ? n10886_o : n10885_o;
  /* TG68K_ALU.vhd:530:30  */
  assign n10888_o = bf_loffset[0];
  /* TG68K_ALU.vhd:531:47  */
  assign n10890_o = {1'b1, bitmaskmux0};
  /* TG68K_ALU.vhd:531:59  */
  assign n10892_o = {n10890_o, 1'b1};
  /* TG68K_ALU.vhd:533:66  */
  assign n10893_o = bitmaskmux0[31];
  assign n10894_o = n10892_o[0];
  /* TG68K_ALU.vhd:532:25  */
  assign n10895_o = bf_d32 ? n10893_o : n10894_o;
  assign n10896_o = n10892_o[39:1];
  /* TG68K_ALU.vhd:536:48  */
  assign n10898_o = {2'b11, bitmaskmux0};
  assign n10899_o = {n10896_o, n10895_o};
  /* TG68K_ALU.vhd:530:17  */
  assign n10900_o = n10888_o ? n10899_o : n10898_o;
  /* TG68K_ALU.vhd:541:35  */
  assign n10901_o = {bf_ext_in, op2out};
  /* TG68K_ALU.vhd:543:54  */
  assign n10902_o = op2out[7:0];
  assign n10903_o = n10901_o[39:32];
  /* TG68K_ALU.vhd:542:17  */
  assign n10904_o = bf_s32 ? n10902_o : n10903_o;
  assign n10905_o = n10901_o[31:0];
  /* TG68K_ALU.vhd:546:28  */
  assign n10906_o = bf_shift[0];
  /* TG68K_ALU.vhd:547:40  */
  assign n10907_o = shift[0];
  /* TG68K_ALU.vhd:547:49  */
  assign n10908_o = shift[39:1];
  /* TG68K_ALU.vhd:547:43  */
  assign n10909_o = {n10907_o, n10908_o};
  /* TG68K_ALU.vhd:546:17  */
  assign n10910_o = n10906_o ? n10909_o : shift;
  /* TG68K_ALU.vhd:551:28  */
  assign n10911_o = bf_shift[1];
  /* TG68K_ALU.vhd:552:41  */
  assign n10912_o = inmux0[1:0];
  /* TG68K_ALU.vhd:552:60  */
  assign n10913_o = inmux0[39:2];
  /* TG68K_ALU.vhd:552:53  */
  assign n10914_o = {n10912_o, n10913_o};
  /* TG68K_ALU.vhd:551:17  */
  assign n10915_o = n10911_o ? n10914_o : inmux0;
  /* TG68K_ALU.vhd:556:28  */
  assign n10916_o = bf_shift[2];
  /* TG68K_ALU.vhd:557:41  */
  assign n10917_o = inmux1[3:0];
  /* TG68K_ALU.vhd:557:60  */
  assign n10918_o = inmux1[39:4];
  /* TG68K_ALU.vhd:557:53  */
  assign n10919_o = {n10917_o, n10918_o};
  /* TG68K_ALU.vhd:556:17  */
  assign n10920_o = n10916_o ? n10919_o : inmux1;
  /* TG68K_ALU.vhd:561:28  */
  assign n10921_o = bf_shift[3];
  /* TG68K_ALU.vhd:562:41  */
  assign n10922_o = inmux2[7:0];
  /* TG68K_ALU.vhd:562:60  */
  assign n10923_o = inmux2[31:8];
  /* TG68K_ALU.vhd:562:53  */
  assign n10924_o = {n10922_o, n10923_o};
  /* TG68K_ALU.vhd:564:41  */
  assign n10925_o = inmux2[31:0];
  /* TG68K_ALU.vhd:561:17  */
  assign n10926_o = n10921_o ? n10924_o : n10925_o;
  /* TG68K_ALU.vhd:566:28  */
  assign n10927_o = bf_shift[4];
  /* TG68K_ALU.vhd:567:55  */
  assign n10928_o = inmux3[15:0];
  /* TG68K_ALU.vhd:567:75  */
  assign n10929_o = inmux3[31:16];
  /* TG68K_ALU.vhd:567:68  */
  assign n10930_o = {n10928_o, n10929_o};
  /* TG68K_ALU.vhd:566:17  */
  assign n10931_o = n10927_o ? n10930_o : inmux3;
  /* TG68K_ALU.vhd:574:56  */
  assign n10932_o = bf_set2[7:0];
  /* TG68K_ALU.vhd:576:48  */
  assign n10933_o = ~op2out;
  /* TG68K_ALU.vhd:577:49  */
  assign n10934_o = ~bf_ext_in;
  assign n10935_o = {n10934_o, n10933_o};
  assign n10938_o = {n10932_o, bf_set2};
  /* TG68K_ALU.vhd:586:48  */
  assign n10942_o = {bf_ext_in, op1out};
  /* TG68K_ALU.vhd:588:48  */
  assign n10943_o = {bf_ext_in, op2out};
  /* TG68K_ALU.vhd:585:17  */
  assign n10944_o = bf_ins ? n10942_o : n10943_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10945_o = shifted_bitmask[0];
  /* TG68K_ALU.vhd:592:56  */
  assign n10946_o = result_tmp[0];
  assign n10947_o = n10940_o[0];
  assign n10948_o = n10938_o[0];
  assign n10949_o = n10935_o[0];
  assign n10950_o = n10936_o[0];
  /* TG68K_ALU.vhd:575:17  */
  assign n10951_o = bf_bchg ? n10949_o : n10950_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10952_o = bf_ins ? n10948_o : n10951_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10953_o = bf_bset ? n10947_o : n10952_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10954_o = n10945_o ? n10946_o : n10953_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10962_o = shifted_bitmask[1];
  /* TG68K_ALU.vhd:592:56  */
  assign n10963_o = result_tmp[1];
  assign n10964_o = n10940_o[1];
  assign n10965_o = n10938_o[1];
  assign n10966_o = n10935_o[1];
  assign n10967_o = n10936_o[1];
  /* TG68K_ALU.vhd:575:17  */
  assign n10968_o = bf_bchg ? n10966_o : n10967_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10969_o = bf_ins ? n10965_o : n10968_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10970_o = bf_bset ? n10964_o : n10969_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10971_o = n10962_o ? n10963_o : n10970_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10979_o = shifted_bitmask[2];
  /* TG68K_ALU.vhd:592:56  */
  assign n10980_o = result_tmp[2];
  assign n10981_o = n10940_o[2];
  assign n10982_o = n10938_o[2];
  assign n10983_o = n10935_o[2];
  assign n10984_o = n10936_o[2];
  /* TG68K_ALU.vhd:575:17  */
  assign n10985_o = bf_bchg ? n10983_o : n10984_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10986_o = bf_ins ? n10982_o : n10985_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10987_o = bf_bset ? n10981_o : n10986_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10988_o = n10979_o ? n10980_o : n10987_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10996_o = shifted_bitmask[3];
  /* TG68K_ALU.vhd:592:56  */
  assign n10997_o = result_tmp[3];
  assign n10998_o = n10940_o[3];
  assign n10999_o = n10938_o[3];
  assign n11000_o = n10935_o[3];
  assign n11001_o = n10936_o[3];
  /* TG68K_ALU.vhd:575:17  */
  assign n11002_o = bf_bchg ? n11000_o : n11001_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11003_o = bf_ins ? n10999_o : n11002_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11004_o = bf_bset ? n10998_o : n11003_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11005_o = n10996_o ? n10997_o : n11004_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11013_o = shifted_bitmask[4];
  /* TG68K_ALU.vhd:592:56  */
  assign n11014_o = result_tmp[4];
  assign n11015_o = n10940_o[4];
  assign n11016_o = n10938_o[4];
  assign n11017_o = n10935_o[4];
  assign n11018_o = n10936_o[4];
  /* TG68K_ALU.vhd:575:17  */
  assign n11019_o = bf_bchg ? n11017_o : n11018_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11020_o = bf_ins ? n11016_o : n11019_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11021_o = bf_bset ? n11015_o : n11020_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11022_o = n11013_o ? n11014_o : n11021_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11030_o = shifted_bitmask[5];
  /* TG68K_ALU.vhd:592:56  */
  assign n11031_o = result_tmp[5];
  assign n11032_o = n10940_o[5];
  assign n11033_o = n10938_o[5];
  assign n11034_o = n10935_o[5];
  assign n11035_o = n10936_o[5];
  /* TG68K_ALU.vhd:575:17  */
  assign n11036_o = bf_bchg ? n11034_o : n11035_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11037_o = bf_ins ? n11033_o : n11036_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11038_o = bf_bset ? n11032_o : n11037_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11039_o = n11030_o ? n11031_o : n11038_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11047_o = shifted_bitmask[6];
  /* TG68K_ALU.vhd:592:56  */
  assign n11048_o = result_tmp[6];
  assign n11049_o = n10940_o[6];
  assign n11050_o = n10938_o[6];
  assign n11051_o = n10935_o[6];
  assign n11052_o = n10936_o[6];
  /* TG68K_ALU.vhd:575:17  */
  assign n11053_o = bf_bchg ? n11051_o : n11052_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11054_o = bf_ins ? n11050_o : n11053_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11055_o = bf_bset ? n11049_o : n11054_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11056_o = n11047_o ? n11048_o : n11055_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11064_o = shifted_bitmask[7];
  /* TG68K_ALU.vhd:592:56  */
  assign n11065_o = result_tmp[7];
  assign n11066_o = n10940_o[7];
  assign n11067_o = n10938_o[7];
  assign n11068_o = n10935_o[7];
  assign n11069_o = n10936_o[7];
  /* TG68K_ALU.vhd:575:17  */
  assign n11070_o = bf_bchg ? n11068_o : n11069_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11071_o = bf_ins ? n11067_o : n11070_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11072_o = bf_bset ? n11066_o : n11071_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11073_o = n11064_o ? n11065_o : n11072_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11081_o = shifted_bitmask[8];
  /* TG68K_ALU.vhd:592:56  */
  assign n11082_o = result_tmp[8];
  assign n11083_o = n10940_o[8];
  assign n11084_o = n10938_o[8];
  assign n11085_o = n10935_o[8];
  assign n11086_o = n10936_o[8];
  /* TG68K_ALU.vhd:575:17  */
  assign n11087_o = bf_bchg ? n11085_o : n11086_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11088_o = bf_ins ? n11084_o : n11087_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11089_o = bf_bset ? n11083_o : n11088_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11090_o = n11081_o ? n11082_o : n11089_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11098_o = shifted_bitmask[9];
  /* TG68K_ALU.vhd:592:56  */
  assign n11099_o = result_tmp[9];
  assign n11100_o = n10940_o[9];
  assign n11101_o = n10938_o[9];
  assign n11102_o = n10935_o[9];
  assign n11103_o = n10936_o[9];
  /* TG68K_ALU.vhd:575:17  */
  assign n11104_o = bf_bchg ? n11102_o : n11103_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11105_o = bf_ins ? n11101_o : n11104_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11106_o = bf_bset ? n11100_o : n11105_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11107_o = n11098_o ? n11099_o : n11106_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11115_o = shifted_bitmask[10];
  /* TG68K_ALU.vhd:592:56  */
  assign n11116_o = result_tmp[10];
  assign n11117_o = n10940_o[10];
  assign n11118_o = n10938_o[10];
  assign n11119_o = n10935_o[10];
  assign n11120_o = n10936_o[10];
  /* TG68K_ALU.vhd:575:17  */
  assign n11121_o = bf_bchg ? n11119_o : n11120_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11122_o = bf_ins ? n11118_o : n11121_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11123_o = bf_bset ? n11117_o : n11122_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11124_o = n11115_o ? n11116_o : n11123_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11132_o = shifted_bitmask[11];
  /* TG68K_ALU.vhd:592:56  */
  assign n11133_o = result_tmp[11];
  assign n11134_o = n10940_o[11];
  assign n11135_o = n10938_o[11];
  assign n11136_o = n10935_o[11];
  assign n11137_o = n10936_o[11];
  /* TG68K_ALU.vhd:575:17  */
  assign n11138_o = bf_bchg ? n11136_o : n11137_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11139_o = bf_ins ? n11135_o : n11138_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11140_o = bf_bset ? n11134_o : n11139_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11141_o = n11132_o ? n11133_o : n11140_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11149_o = shifted_bitmask[12];
  /* TG68K_ALU.vhd:592:56  */
  assign n11150_o = result_tmp[12];
  assign n11151_o = n10940_o[12];
  assign n11152_o = n10938_o[12];
  assign n11153_o = n10935_o[12];
  assign n11154_o = n10936_o[12];
  /* TG68K_ALU.vhd:575:17  */
  assign n11155_o = bf_bchg ? n11153_o : n11154_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11156_o = bf_ins ? n11152_o : n11155_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11157_o = bf_bset ? n11151_o : n11156_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11158_o = n11149_o ? n11150_o : n11157_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11166_o = shifted_bitmask[13];
  /* TG68K_ALU.vhd:592:56  */
  assign n11167_o = result_tmp[13];
  assign n11168_o = n10940_o[13];
  assign n11169_o = n10938_o[13];
  assign n11170_o = n10935_o[13];
  assign n11171_o = n10936_o[13];
  /* TG68K_ALU.vhd:575:17  */
  assign n11172_o = bf_bchg ? n11170_o : n11171_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11173_o = bf_ins ? n11169_o : n11172_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11174_o = bf_bset ? n11168_o : n11173_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11175_o = n11166_o ? n11167_o : n11174_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11183_o = shifted_bitmask[14];
  /* TG68K_ALU.vhd:592:56  */
  assign n11184_o = result_tmp[14];
  assign n11185_o = n10940_o[14];
  assign n11186_o = n10938_o[14];
  assign n11187_o = n10935_o[14];
  assign n11188_o = n10936_o[14];
  /* TG68K_ALU.vhd:575:17  */
  assign n11189_o = bf_bchg ? n11187_o : n11188_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11190_o = bf_ins ? n11186_o : n11189_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11191_o = bf_bset ? n11185_o : n11190_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11192_o = n11183_o ? n11184_o : n11191_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11200_o = shifted_bitmask[15];
  /* TG68K_ALU.vhd:592:56  */
  assign n11201_o = result_tmp[15];
  assign n11202_o = n10940_o[15];
  assign n11203_o = n10938_o[15];
  assign n11204_o = n10935_o[15];
  assign n11205_o = n10936_o[15];
  /* TG68K_ALU.vhd:575:17  */
  assign n11206_o = bf_bchg ? n11204_o : n11205_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11207_o = bf_ins ? n11203_o : n11206_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11208_o = bf_bset ? n11202_o : n11207_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11209_o = n11200_o ? n11201_o : n11208_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11217_o = shifted_bitmask[16];
  /* TG68K_ALU.vhd:592:56  */
  assign n11218_o = result_tmp[16];
  assign n11219_o = n10940_o[16];
  assign n11220_o = n10938_o[16];
  assign n11221_o = n10935_o[16];
  assign n11222_o = n10936_o[16];
  /* TG68K_ALU.vhd:575:17  */
  assign n11223_o = bf_bchg ? n11221_o : n11222_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11224_o = bf_ins ? n11220_o : n11223_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11225_o = bf_bset ? n11219_o : n11224_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11226_o = n11217_o ? n11218_o : n11225_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11234_o = shifted_bitmask[17];
  /* TG68K_ALU.vhd:592:56  */
  assign n11235_o = result_tmp[17];
  assign n11236_o = n10940_o[17];
  assign n11237_o = n10938_o[17];
  assign n11238_o = n10935_o[17];
  assign n11239_o = n10936_o[17];
  /* TG68K_ALU.vhd:575:17  */
  assign n11240_o = bf_bchg ? n11238_o : n11239_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11241_o = bf_ins ? n11237_o : n11240_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11242_o = bf_bset ? n11236_o : n11241_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11243_o = n11234_o ? n11235_o : n11242_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11251_o = shifted_bitmask[18];
  /* TG68K_ALU.vhd:592:56  */
  assign n11252_o = result_tmp[18];
  assign n11253_o = n10940_o[18];
  assign n11254_o = n10938_o[18];
  assign n11255_o = n10935_o[18];
  assign n11256_o = n10936_o[18];
  /* TG68K_ALU.vhd:575:17  */
  assign n11257_o = bf_bchg ? n11255_o : n11256_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11258_o = bf_ins ? n11254_o : n11257_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11259_o = bf_bset ? n11253_o : n11258_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11260_o = n11251_o ? n11252_o : n11259_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11268_o = shifted_bitmask[19];
  /* TG68K_ALU.vhd:592:56  */
  assign n11269_o = result_tmp[19];
  assign n11270_o = n10940_o[19];
  assign n11271_o = n10938_o[19];
  assign n11272_o = n10935_o[19];
  assign n11273_o = n10936_o[19];
  /* TG68K_ALU.vhd:575:17  */
  assign n11274_o = bf_bchg ? n11272_o : n11273_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11275_o = bf_ins ? n11271_o : n11274_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11276_o = bf_bset ? n11270_o : n11275_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11277_o = n11268_o ? n11269_o : n11276_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11285_o = shifted_bitmask[20];
  /* TG68K_ALU.vhd:592:56  */
  assign n11286_o = result_tmp[20];
  assign n11287_o = n10940_o[20];
  assign n11288_o = n10938_o[20];
  assign n11289_o = n10935_o[20];
  assign n11290_o = n10936_o[20];
  /* TG68K_ALU.vhd:575:17  */
  assign n11291_o = bf_bchg ? n11289_o : n11290_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11292_o = bf_ins ? n11288_o : n11291_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11293_o = bf_bset ? n11287_o : n11292_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11294_o = n11285_o ? n11286_o : n11293_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11302_o = shifted_bitmask[21];
  /* TG68K_ALU.vhd:592:56  */
  assign n11303_o = result_tmp[21];
  assign n11304_o = n10940_o[21];
  assign n11305_o = n10938_o[21];
  assign n11306_o = n10935_o[21];
  assign n11307_o = n10936_o[21];
  /* TG68K_ALU.vhd:575:17  */
  assign n11308_o = bf_bchg ? n11306_o : n11307_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11309_o = bf_ins ? n11305_o : n11308_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11310_o = bf_bset ? n11304_o : n11309_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11311_o = n11302_o ? n11303_o : n11310_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11319_o = shifted_bitmask[22];
  /* TG68K_ALU.vhd:592:56  */
  assign n11320_o = result_tmp[22];
  assign n11321_o = n10940_o[22];
  assign n11322_o = n10938_o[22];
  assign n11323_o = n10935_o[22];
  assign n11324_o = n10936_o[22];
  /* TG68K_ALU.vhd:575:17  */
  assign n11325_o = bf_bchg ? n11323_o : n11324_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11326_o = bf_ins ? n11322_o : n11325_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11327_o = bf_bset ? n11321_o : n11326_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11328_o = n11319_o ? n11320_o : n11327_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11336_o = shifted_bitmask[23];
  /* TG68K_ALU.vhd:592:56  */
  assign n11337_o = result_tmp[23];
  assign n11338_o = n10940_o[23];
  assign n11339_o = n10938_o[23];
  assign n11340_o = n10935_o[23];
  assign n11341_o = n10936_o[23];
  /* TG68K_ALU.vhd:575:17  */
  assign n11342_o = bf_bchg ? n11340_o : n11341_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11343_o = bf_ins ? n11339_o : n11342_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11344_o = bf_bset ? n11338_o : n11343_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11345_o = n11336_o ? n11337_o : n11344_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11353_o = shifted_bitmask[24];
  /* TG68K_ALU.vhd:592:56  */
  assign n11354_o = result_tmp[24];
  assign n11355_o = n10940_o[24];
  assign n11356_o = n10938_o[24];
  assign n11357_o = n10935_o[24];
  assign n11358_o = n10936_o[24];
  /* TG68K_ALU.vhd:575:17  */
  assign n11359_o = bf_bchg ? n11357_o : n11358_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11360_o = bf_ins ? n11356_o : n11359_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11361_o = bf_bset ? n11355_o : n11360_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11362_o = n11353_o ? n11354_o : n11361_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11370_o = shifted_bitmask[25];
  /* TG68K_ALU.vhd:592:56  */
  assign n11371_o = result_tmp[25];
  assign n11372_o = n10940_o[25];
  assign n11373_o = n10938_o[25];
  assign n11374_o = n10935_o[25];
  assign n11375_o = n10936_o[25];
  /* TG68K_ALU.vhd:575:17  */
  assign n11376_o = bf_bchg ? n11374_o : n11375_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11377_o = bf_ins ? n11373_o : n11376_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11378_o = bf_bset ? n11372_o : n11377_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11379_o = n11370_o ? n11371_o : n11378_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11387_o = shifted_bitmask[26];
  /* TG68K_ALU.vhd:592:56  */
  assign n11388_o = result_tmp[26];
  assign n11389_o = n10940_o[26];
  assign n11390_o = n10938_o[26];
  assign n11391_o = n10935_o[26];
  assign n11392_o = n10936_o[26];
  /* TG68K_ALU.vhd:575:17  */
  assign n11393_o = bf_bchg ? n11391_o : n11392_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11394_o = bf_ins ? n11390_o : n11393_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11395_o = bf_bset ? n11389_o : n11394_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11396_o = n11387_o ? n11388_o : n11395_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11404_o = shifted_bitmask[27];
  /* TG68K_ALU.vhd:592:56  */
  assign n11405_o = result_tmp[27];
  assign n11406_o = n10940_o[27];
  assign n11407_o = n10938_o[27];
  assign n11408_o = n10935_o[27];
  assign n11409_o = n10936_o[27];
  /* TG68K_ALU.vhd:575:17  */
  assign n11410_o = bf_bchg ? n11408_o : n11409_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11411_o = bf_ins ? n11407_o : n11410_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11412_o = bf_bset ? n11406_o : n11411_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11413_o = n11404_o ? n11405_o : n11412_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11421_o = shifted_bitmask[28];
  /* TG68K_ALU.vhd:592:56  */
  assign n11422_o = result_tmp[28];
  assign n11423_o = n10940_o[28];
  assign n11424_o = n10938_o[28];
  assign n11425_o = n10935_o[28];
  assign n11426_o = n10936_o[28];
  /* TG68K_ALU.vhd:575:17  */
  assign n11427_o = bf_bchg ? n11425_o : n11426_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11428_o = bf_ins ? n11424_o : n11427_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11429_o = bf_bset ? n11423_o : n11428_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11430_o = n11421_o ? n11422_o : n11429_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11438_o = shifted_bitmask[29];
  /* TG68K_ALU.vhd:592:56  */
  assign n11439_o = result_tmp[29];
  assign n11440_o = n10940_o[29];
  assign n11441_o = n10938_o[29];
  assign n11442_o = n10935_o[29];
  assign n11443_o = n10936_o[29];
  /* TG68K_ALU.vhd:575:17  */
  assign n11444_o = bf_bchg ? n11442_o : n11443_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11445_o = bf_ins ? n11441_o : n11444_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11446_o = bf_bset ? n11440_o : n11445_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11447_o = n11438_o ? n11439_o : n11446_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11455_o = shifted_bitmask[30];
  /* TG68K_ALU.vhd:592:56  */
  assign n11456_o = result_tmp[30];
  assign n11457_o = n10940_o[30];
  assign n11458_o = n10938_o[30];
  assign n11459_o = n10935_o[30];
  assign n11460_o = n10936_o[30];
  /* TG68K_ALU.vhd:575:17  */
  assign n11461_o = bf_bchg ? n11459_o : n11460_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11462_o = bf_ins ? n11458_o : n11461_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11463_o = bf_bset ? n11457_o : n11462_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11464_o = n11455_o ? n11456_o : n11463_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11472_o = shifted_bitmask[31];
  /* TG68K_ALU.vhd:592:56  */
  assign n11473_o = result_tmp[31];
  assign n11474_o = n10940_o[31];
  assign n11475_o = n10938_o[31];
  assign n11476_o = n10935_o[31];
  assign n11477_o = n10936_o[31];
  /* TG68K_ALU.vhd:575:17  */
  assign n11478_o = bf_bchg ? n11476_o : n11477_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11479_o = bf_ins ? n11475_o : n11478_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11480_o = bf_bset ? n11474_o : n11479_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11481_o = n11472_o ? n11473_o : n11480_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11489_o = shifted_bitmask[32];
  /* TG68K_ALU.vhd:592:56  */
  assign n11490_o = result_tmp[32];
  assign n11491_o = n10940_o[32];
  assign n11492_o = n10938_o[32];
  assign n11493_o = n10935_o[32];
  assign n11494_o = n10936_o[32];
  /* TG68K_ALU.vhd:575:17  */
  assign n11495_o = bf_bchg ? n11493_o : n11494_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11496_o = bf_ins ? n11492_o : n11495_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11497_o = bf_bset ? n11491_o : n11496_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11498_o = n11489_o ? n11490_o : n11497_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11506_o = shifted_bitmask[33];
  /* TG68K_ALU.vhd:592:56  */
  assign n11507_o = result_tmp[33];
  assign n11508_o = n10940_o[33];
  assign n11509_o = n10938_o[33];
  assign n11510_o = n10935_o[33];
  assign n11511_o = n10936_o[33];
  /* TG68K_ALU.vhd:575:17  */
  assign n11512_o = bf_bchg ? n11510_o : n11511_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11513_o = bf_ins ? n11509_o : n11512_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11514_o = bf_bset ? n11508_o : n11513_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11515_o = n11506_o ? n11507_o : n11514_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11523_o = shifted_bitmask[34];
  /* TG68K_ALU.vhd:592:56  */
  assign n11524_o = result_tmp[34];
  assign n11525_o = n10940_o[34];
  assign n11526_o = n10938_o[34];
  assign n11527_o = n10935_o[34];
  assign n11528_o = n10936_o[34];
  /* TG68K_ALU.vhd:575:17  */
  assign n11529_o = bf_bchg ? n11527_o : n11528_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11530_o = bf_ins ? n11526_o : n11529_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11531_o = bf_bset ? n11525_o : n11530_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11532_o = n11523_o ? n11524_o : n11531_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11540_o = shifted_bitmask[35];
  /* TG68K_ALU.vhd:592:56  */
  assign n11541_o = result_tmp[35];
  assign n11542_o = n10940_o[35];
  assign n11543_o = n10938_o[35];
  assign n11544_o = n10935_o[35];
  assign n11545_o = n10936_o[35];
  /* TG68K_ALU.vhd:575:17  */
  assign n11546_o = bf_bchg ? n11544_o : n11545_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11547_o = bf_ins ? n11543_o : n11546_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11548_o = bf_bset ? n11542_o : n11547_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11549_o = n11540_o ? n11541_o : n11548_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11557_o = shifted_bitmask[36];
  /* TG68K_ALU.vhd:592:56  */
  assign n11558_o = result_tmp[36];
  assign n11559_o = n10940_o[36];
  assign n11560_o = n10938_o[36];
  assign n11561_o = n10935_o[36];
  assign n11562_o = n10936_o[36];
  /* TG68K_ALU.vhd:575:17  */
  assign n11563_o = bf_bchg ? n11561_o : n11562_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11564_o = bf_ins ? n11560_o : n11563_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11565_o = bf_bset ? n11559_o : n11564_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11566_o = n11557_o ? n11558_o : n11565_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11574_o = shifted_bitmask[37];
  /* TG68K_ALU.vhd:592:56  */
  assign n11575_o = result_tmp[37];
  assign n11576_o = n10940_o[37];
  assign n11577_o = n10938_o[37];
  assign n11578_o = n10935_o[37];
  assign n11579_o = n10936_o[37];
  /* TG68K_ALU.vhd:575:17  */
  assign n11580_o = bf_bchg ? n11578_o : n11579_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11581_o = bf_ins ? n11577_o : n11580_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11582_o = bf_bset ? n11576_o : n11581_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11583_o = n11574_o ? n11575_o : n11582_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11591_o = shifted_bitmask[38];
  /* TG68K_ALU.vhd:592:56  */
  assign n11592_o = result_tmp[38];
  assign n11593_o = n10940_o[38];
  assign n11594_o = n10938_o[38];
  assign n11595_o = n10935_o[38];
  assign n11596_o = n10936_o[38];
  /* TG68K_ALU.vhd:575:17  */
  assign n11597_o = bf_bchg ? n11595_o : n11596_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11598_o = bf_ins ? n11594_o : n11597_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11599_o = bf_bset ? n11593_o : n11598_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11600_o = n11591_o ? n11592_o : n11599_o;
  assign n11601_o = n10940_o[39];
  assign n11602_o = n10938_o[39];
  assign n11603_o = n10935_o[39];
  assign n11604_o = n10936_o[39];
  /* TG68K_ALU.vhd:575:17  */
  assign n11605_o = bf_bchg ? n11603_o : n11604_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11606_o = bf_ins ? n11602_o : n11605_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11607_o = bf_bset ? n11601_o : n11606_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11608_o = shifted_bitmask[39];
  /* TG68K_ALU.vhd:592:56  */
  assign n11609_o = result_tmp[39];
  /* TG68K_ALU.vhd:591:25  */
  assign n11610_o = n11608_o ? n11609_o : n11607_o;
  /* TG68K_ALU.vhd:598:36  */
  assign n11612_o = {1'b0, bitnr};
  /* TG68K_ALU.vhd:598:43  */
  assign n11613_o = {5'b0, mask_not_zero};  //  uext
  /* TG68K_ALU.vhd:598:43  */
  assign n11614_o = n11612_o + n11613_o;
  /* TG68K_ALU.vhd:601:24  */
  assign n11615_o = mask[31:28];
  /* TG68K_ALU.vhd:601:38  */
  assign n11617_o = n11615_o == 4'b0000;
  /* TG68K_ALU.vhd:602:32  */
  assign n11618_o = mask[27:24];
  /* TG68K_ALU.vhd:602:46  */
  assign n11620_o = n11618_o == 4'b0000;
  /* TG68K_ALU.vhd:603:40  */
  assign n11621_o = mask[23:20];
  /* TG68K_ALU.vhd:603:54  */
  assign n11623_o = n11621_o == 4'b0000;
  /* TG68K_ALU.vhd:604:48  */
  assign n11624_o = mask[19:16];
  /* TG68K_ALU.vhd:604:62  */
  assign n11626_o = n11624_o == 4'b0000;
  /* TG68K_ALU.vhd:606:56  */
  assign n11628_o = mask[15:12];
  /* TG68K_ALU.vhd:606:70  */
  assign n11630_o = n11628_o == 4'b0000;
  /* TG68K_ALU.vhd:607:64  */
  assign n11631_o = mask[11:8];
  /* TG68K_ALU.vhd:607:77  */
  assign n11633_o = n11631_o == 4'b0000;
  /* TG68K_ALU.vhd:609:72  */
  assign n11635_o = mask[7:4];
  /* TG68K_ALU.vhd:609:84  */
  assign n11637_o = n11635_o == 4'b0000;
  /* TG68K_ALU.vhd:611:84  */
  assign n11639_o = mask[3:0];
  /* TG68K_ALU.vhd:613:84  */
  assign n11640_o = mask[7:4];
  /* TG68K_ALU.vhd:609:65  */
  assign n11641_o = n11637_o ? n11639_o : n11640_o;
  /* TG68K_ALU.vhd:609:65  */
  assign n11643_o = n11637_o ? 1'b0 : 1'b1;
  /* TG68K_ALU.vhd:616:76  */
  assign n11644_o = mask[11:8];
  /* TG68K_ALU.vhd:607:57  */
  assign n11646_o = n11633_o ? n11641_o : n11644_o;
  assign n11647_o = {1'b0, n11643_o};
  assign n11648_o = n11647_o[0];
  /* TG68K_ALU.vhd:607:57  */
  assign n11649_o = n11633_o ? n11648_o : 1'b0;
  assign n11650_o = n11647_o[1];
  /* TG68K_ALU.vhd:607:57  */
  assign n11652_o = n11633_o ? n11650_o : 1'b1;
  /* TG68K_ALU.vhd:620:68  */
  assign n11653_o = mask[15:12];
  /* TG68K_ALU.vhd:606:49  */
  assign n11654_o = n11630_o ? n11646_o : n11653_o;
  assign n11655_o = {n11652_o, n11649_o};
  /* TG68K_ALU.vhd:606:49  */
  assign n11657_o = n11630_o ? n11655_o : 2'b11;
  /* TG68K_ALU.vhd:623:60  */
  assign n11658_o = mask[19:16];
  /* TG68K_ALU.vhd:604:41  */
  assign n11661_o = n11626_o ? n11654_o : n11658_o;
  assign n11662_o = {1'b0, 1'b0};
  assign n11663_o = {1'b0, n11657_o};
  assign n11664_o = n11663_o[1:0];
  /* TG68K_ALU.vhd:604:41  */
  assign n11665_o = n11626_o ? n11664_o : n11662_o;
  assign n11666_o = n11663_o[2];
  /* TG68K_ALU.vhd:604:41  */
  assign n11668_o = n11626_o ? n11666_o : 1'b1;
  /* TG68K_ALU.vhd:628:52  */
  assign n11669_o = mask[23:20];
  /* TG68K_ALU.vhd:603:33  */
  assign n11671_o = n11623_o ? n11661_o : n11669_o;
  assign n11672_o = {n11668_o, n11665_o};
  assign n11673_o = n11672_o[0];
  /* TG68K_ALU.vhd:603:33  */
  assign n11675_o = n11623_o ? n11673_o : 1'b1;
  assign n11676_o = n11672_o[1];
  /* TG68K_ALU.vhd:603:33  */
  assign n11677_o = n11623_o ? n11676_o : 1'b0;
  assign n11678_o = n11672_o[2];
  /* TG68K_ALU.vhd:603:33  */
  assign n11680_o = n11623_o ? n11678_o : 1'b1;
  /* TG68K_ALU.vhd:632:44  */
  assign n11681_o = mask[27:24];
  /* TG68K_ALU.vhd:602:25  */
  assign n11683_o = n11620_o ? n11671_o : n11681_o;
  assign n11684_o = {n11680_o, n11677_o, n11675_o};
  assign n11685_o = n11684_o[0];
  /* TG68K_ALU.vhd:602:25  */
  assign n11686_o = n11620_o ? n11685_o : 1'b0;
  assign n11687_o = n11684_o[2:1];
  /* TG68K_ALU.vhd:602:25  */
  assign n11689_o = n11620_o ? n11687_o : 2'b11;
  /* TG68K_ALU.vhd:636:36  */
  assign n11690_o = mask[31:28];
  /* TG68K_ALU.vhd:601:17  */
  assign n11691_o = n11617_o ? n11683_o : n11690_o;
  assign n11692_o = {n11689_o, n11686_o};
  /* TG68K_ALU.vhd:601:17  */
  assign n11694_o = n11617_o ? n11692_o : 3'b111;
  /* TG68K_ALU.vhd:639:23  */
  assign n11697_o = mux[3:2];
  /* TG68K_ALU.vhd:639:35  */
  assign n11699_o = n11697_o == 2'b00;
  /* TG68K_ALU.vhd:641:31  */
  assign n11701_o = mux[1];
  /* TG68K_ALU.vhd:641:34  */
  assign n11702_o = ~n11701_o;
  /* TG68K_ALU.vhd:643:39  */
  assign n11704_o = mux[0];
  /* TG68K_ALU.vhd:643:42  */
  assign n11705_o = ~n11704_o;
  /* TG68K_ALU.vhd:643:33  */
  assign n11708_o = n11705_o ? 1'b0 : 1'b1;
  assign n11709_o = n11695_o[0];
  /* TG68K_ALU.vhd:641:25  */
  assign n11710_o = n11702_o ? 1'b0 : n11709_o;
  /* TG68K_ALU.vhd:641:25  */
  assign n11712_o = n11702_o ? n11708_o : 1'b1;
  /* TG68K_ALU.vhd:648:31  */
  assign n11713_o = mux[3];
  /* TG68K_ALU.vhd:648:34  */
  assign n11714_o = ~n11713_o;
  assign n11716_o = n11695_o[0];
  /* TG68K_ALU.vhd:648:25  */
  assign n11717_o = n11714_o ? 1'b0 : n11716_o;
  assign n11718_o = {1'b0, n11710_o};
  assign n11719_o = n11718_o[0];
  /* TG68K_ALU.vhd:639:17  */
  assign n11720_o = n11699_o ? n11719_o : n11717_o;
  assign n11721_o = n11718_o[1];
  assign n11722_o = n11695_o[1];
  /* TG68K_ALU.vhd:639:17  */
  assign n11723_o = n11699_o ? n11721_o : n11722_o;
  /* TG68K_ALU.vhd:639:17  */
  assign n11726_o = n11699_o ? n11712_o : 1'b1;
  /* TG68K_ALU.vhd:659:32  */
  assign n11731_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:661:66  */
  assign n11732_o = op1out[7];
  /* TG68K_ALU.vhd:660:25  */
  assign n11734_o = n11731_o == 2'b00;
  /* TG68K_ALU.vhd:663:66  */
  assign n11735_o = op1out[15];
  /* TG68K_ALU.vhd:662:25  */
  assign n11737_o = n11731_o == 2'b01;
  /* TG68K_ALU.vhd:662:34  */
  assign n11739_o = n11731_o == 2'b11;
  /* TG68K_ALU.vhd:662:34  */
  assign n11740_o = n11737_o | n11739_o;
  /* TG68K_ALU.vhd:665:66  */
  assign n11741_o = op1out[31];
  /* TG68K_ALU.vhd:664:25  */
  assign n11743_o = n11731_o == 2'b10;
  assign n11744_o = {n11743_o, n11740_o, n11734_o};
  /* TG68K_ALU.vhd:659:17  */
  always @*
    case (n11744_o)
      3'b100: n11745_o = n11741_o;
      3'b010: n11745_o = n11735_o;
      3'b001: n11745_o = n11732_o;
      default: n11745_o = rot_rot;
    endcase
  /* TG68K_ALU.vhd:685:24  */
  assign n11763_o = exec[23];
  /* TG68K_ALU.vhd:687:39  */
  assign n11764_o = n12945_q[4];
  /* TG68K_ALU.vhd:688:36  */
  assign n11766_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:689:47  */
  assign n11767_o = n12945_q[4];
  /* TG68K_ALU.vhd:688:25  */
  assign n11769_o = n11766_o ? n11767_o : 1'b0;
  /* TG68K_ALU.vhd:694:38  */
  assign n11770_o = exe_opcode[8];
  /* TG68K_ALU.vhd:699:48  */
  assign n11773_o = op1out[0];
  /* TG68K_ALU.vhd:700:48  */
  assign n11774_o = op1out[0];
  /* TG68K_ALU.vhd:694:25  */
  assign n11794_o = n11770_o ? rot_rot : n11773_o;
  /* TG68K_ALU.vhd:694:25  */
  assign n11795_o = n11770_o ? rot_rot : n11774_o;
  /* TG68K_ALU.vhd:685:17  */
  assign n11798_o = n11763_o ? n11764_o : n11794_o;
  /* TG68K_ALU.vhd:685:17  */
  assign n11799_o = n11763_o ? n11769_o : n11795_o;
  /* TG68K_ALU.vhd:685:17  */
  assign n11800_o = n11763_o ? op1out : bsout;
  /* TG68K_ALU.vhd:723:28  */
  assign n11805_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:724:40  */
  assign n11806_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:725:33  */
  assign n11808_o = n11806_o == 2'b00;
  /* TG68K_ALU.vhd:727:33  */
  assign n11810_o = n11806_o == 2'b01;
  /* TG68K_ALU.vhd:727:42  */
  assign n11812_o = n11806_o == 2'b11;
  /* TG68K_ALU.vhd:727:42  */
  assign n11813_o = n11810_o | n11812_o;
  /* TG68K_ALU.vhd:729:33  */
  assign n11815_o = n11806_o == 2'b10;
  assign n11816_o = {n11815_o, n11813_o, n11808_o};
  /* TG68K_ALU.vhd:724:25  */
  always @*
    case (n11816_o)
      3'b100: n11821_o = 6'b100001;
      3'b010: n11821_o = 6'b010001;
      3'b001: n11821_o = 6'b001001;
      default: n11821_o = 6'b100000;
    endcase
  /* TG68K_ALU.vhd:734:40  */
  assign n11822_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:735:33  */
  assign n11824_o = n11822_o == 2'b00;
  /* TG68K_ALU.vhd:737:33  */
  assign n11826_o = n11822_o == 2'b01;
  /* TG68K_ALU.vhd:737:42  */
  assign n11828_o = n11822_o == 2'b11;
  /* TG68K_ALU.vhd:737:42  */
  assign n11829_o = n11826_o | n11828_o;
  /* TG68K_ALU.vhd:739:33  */
  assign n11831_o = n11822_o == 2'b10;
  assign n11832_o = {n11831_o, n11829_o, n11824_o};
  /* TG68K_ALU.vhd:734:25  */
  always @*
    case (n11832_o)
      3'b100: n11837_o = 6'b100000;
      3'b010: n11837_o = 6'b010000;
      3'b001: n11837_o = 6'b001000;
      default: n11837_o = 6'b100000;
    endcase
  /* TG68K_ALU.vhd:723:17  */
  assign n11838_o = n11805_o ? n11821_o : n11837_o;
  /* TG68K_ALU.vhd:745:30  */
  assign n11840_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:745:42  */
  assign n11842_o = n11840_o == 2'b11;
  /* TG68K_ALU.vhd:745:55  */
  assign n11843_o = exec[81];
  /* TG68K_ALU.vhd:745:64  */
  assign n11844_o = ~n11843_o;
  /* TG68K_ALU.vhd:745:48  */
  assign n11845_o = n11842_o | n11844_o;
  /* TG68K_ALU.vhd:747:33  */
  assign n11846_o = exe_opcode[5];
  /* TG68K_ALU.vhd:748:43  */
  assign n11847_o = op2out[5:0];
  /* TG68K_ALU.vhd:750:59  */
  assign n11848_o = exe_opcode[11:9];
  /* TG68K_ALU.vhd:751:38  */
  assign n11849_o = exe_opcode[11:9];
  /* TG68K_ALU.vhd:751:51  */
  assign n11851_o = n11849_o == 3'b000;
  /* TG68K_ALU.vhd:751:25  */
  assign n11854_o = n11851_o ? 3'b001 : 3'b000;
  assign n11855_o = {n11854_o, n11848_o};
  /* TG68K_ALU.vhd:747:17  */
  assign n11856_o = n11846_o ? n11847_o : n11855_o;
  /* TG68K_ALU.vhd:745:17  */
  assign n11858_o = n11845_o ? 6'b000001 : n11856_o;
  /* TG68K_ALU.vhd:762:29  */
  assign n11865_o = $unsigned(bs_shift) < $unsigned(ring);
  /* TG68K_ALU.vhd:763:40  */
  assign n11866_o = ring - bs_shift;
  /* TG68K_ALU.vhd:762:17  */
  assign n11868_o = n11865_o ? n11866_o : 6'b000000;
  /* TG68K_ALU.vhd:765:45  */
  assign n11870_o = vector[30:0];
  /* TG68K_ALU.vhd:765:38  */
  assign n11872_o = {1'b0, n11870_o};
  /* TG68K_ALU.vhd:765:75  */
  assign n11873_o = vector[31:1];
  /* TG68K_ALU.vhd:765:68  */
  assign n11875_o = {1'b0, n11873_o};
  /* TG68K_ALU.vhd:765:60  */
  assign n11876_o = n11872_o ^ n11875_o;
  /* TG68K_ALU.vhd:765:90  */
  assign n11877_o = {n11876_o, msb};
  /* TG68K_ALU.vhd:766:32  */
  assign n11878_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:767:25  */
  assign n11881_o = n11878_o == 2'b00;
  /* TG68K_ALU.vhd:769:25  */
  assign n11884_o = n11878_o == 2'b01;
  /* TG68K_ALU.vhd:769:34  */
  assign n11886_o = n11878_o == 2'b11;
  /* TG68K_ALU.vhd:769:34  */
  assign n11887_o = n11884_o | n11886_o;
  assign n11888_o = {n11887_o, n11881_o};
  assign n11889_o = n11877_o[8];
  /* TG68K_ALU.vhd:766:17  */
  always @*
    case (n11888_o)
      2'b10: n11890_o = n11889_o;
      2'b01: n11890_o = 1'b0;
      default: n11890_o = n11889_o;
    endcase
  assign n11891_o = n11877_o[16];
  /* TG68K_ALU.vhd:766:17  */
  always @*
    case (n11888_o)
      2'b10: n11892_o = 1'b0;
      2'b01: n11892_o = n11891_o;
      default: n11892_o = n11891_o;
    endcase
  assign n11894_o = n11877_o[7:0];
  assign n11895_o = n11877_o[32:17];
  assign n11896_o = n11877_o[15:9];
  /* TG68K_ALU.vhd:773:56  */
  assign n11897_o = hot_msb[31:0];
  /* TG68K_ALU.vhd:773:48  */
  assign n11899_o = {1'b0, n11897_o};
  /* TG68K_ALU.vhd:773:42  */
  assign n11900_o = asl_over_xor - n11899_o;
  /* TG68K_ALU.vhd:775:28  */
  assign n11902_o = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:775:48  */
  assign n11903_o = exe_opcode[8];
  /* TG68K_ALU.vhd:775:34  */
  assign n11904_o = n11903_o & n11902_o;
  /* TG68K_ALU.vhd:776:45  */
  assign n11905_o = asl_over[32];
  /* TG68K_ALU.vhd:776:33  */
  assign n11906_o = ~n11905_o;
  /* TG68K_ALU.vhd:775:17  */
  assign n11908_o = n11904_o ? n11906_o : 1'b0;
  /* TG68K_ALU.vhd:780:30  */
  assign n11910_o = exe_opcode[8];
  /* TG68K_ALU.vhd:780:33  */
  assign n11911_o = ~n11910_o;
  /* TG68K_ALU.vhd:781:42  */
  assign n11912_o = result_bs[31];
  /* TG68K_ALU.vhd:783:40  */
  assign n11913_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:785:58  */
  assign n11914_o = result_bs[8];
  /* TG68K_ALU.vhd:784:33  */
  assign n11916_o = n11913_o == 2'b00;
  /* TG68K_ALU.vhd:787:58  */
  assign n11917_o = result_bs[16];
  /* TG68K_ALU.vhd:786:33  */
  assign n11919_o = n11913_o == 2'b01;
  /* TG68K_ALU.vhd:786:42  */
  assign n11921_o = n11913_o == 2'b11;
  /* TG68K_ALU.vhd:786:42  */
  assign n11922_o = n11919_o | n11921_o;
  /* TG68K_ALU.vhd:789:58  */
  assign n11923_o = result_bs[32];
  /* TG68K_ALU.vhd:788:33  */
  assign n11925_o = n11913_o == 2'b10;
  assign n11926_o = {n11925_o, n11922_o, n11916_o};
  /* TG68K_ALU.vhd:783:25  */
  always @*
    case (n11926_o)
      3'b100: n11927_o = n11923_o;
      3'b010: n11927_o = n11917_o;
      3'b001: n11927_o = n11914_o;
      default: n11927_o = bs_c;
    endcase
  /* TG68K_ALU.vhd:780:17  */
  assign n11928_o = n11911_o ? n11912_o : n11927_o;
  /* TG68K_ALU.vhd:795:28  */
  assign n11930_o = rot_bits == 2'b11;
  /* TG68K_ALU.vhd:796:38  */
  assign n11931_o = n12945_q[4];
  /* TG68K_ALU.vhd:797:40  */
  assign n11932_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:799:69  */
  assign n11933_o = result_bs[7:0];
  /* TG68K_ALU.vhd:799:94  */
  assign n11934_o = result_bs[15:8];
  /* TG68K_ALU.vhd:799:82  */
  assign n11935_o = n11933_o | n11934_o;
  /* TG68K_ALU.vhd:800:52  */
  assign n11936_o = alu[7];
  /* TG68K_ALU.vhd:798:33  */
  assign n11938_o = n11932_o == 2'b00;
  /* TG68K_ALU.vhd:802:70  */
  assign n11939_o = result_bs[15:0];
  /* TG68K_ALU.vhd:802:96  */
  assign n11940_o = result_bs[31:16];
  /* TG68K_ALU.vhd:802:84  */
  assign n11941_o = n11939_o | n11940_o;
  /* TG68K_ALU.vhd:803:52  */
  assign n11942_o = alu[15];
  /* TG68K_ALU.vhd:801:33  */
  assign n11944_o = n11932_o == 2'b01;
  /* TG68K_ALU.vhd:801:42  */
  assign n11946_o = n11932_o == 2'b11;
  /* TG68K_ALU.vhd:801:42  */
  assign n11947_o = n11944_o | n11946_o;
  /* TG68K_ALU.vhd:805:57  */
  assign n11948_o = result_bs[31:0];
  /* TG68K_ALU.vhd:805:83  */
  assign n11949_o = result_bs[63:32];
  /* TG68K_ALU.vhd:805:71  */
  assign n11950_o = n11948_o | n11949_o;
  /* TG68K_ALU.vhd:806:52  */
  assign n11951_o = alu[31];
  /* TG68K_ALU.vhd:804:33  */
  assign n11953_o = n11932_o == 2'b10;
  assign n11954_o = {n11953_o, n11947_o, n11938_o};
  assign n11955_o = n11941_o[7:0];
  assign n11956_o = n11950_o[7:0];
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11954_o)
      3'b100: n11958_o = n11956_o;
      3'b010: n11958_o = n11955_o;
      3'b001: n11958_o = n11935_o;
      default: n11958_o = 8'bX;
    endcase
  assign n11959_o = n11941_o[15:8];
  assign n11960_o = n11950_o[15:8];
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11954_o)
      3'b100: n11962_o = n11960_o;
      3'b010: n11962_o = n11959_o;
      3'b001: n11962_o = 8'bX;
      default: n11962_o = 8'bX;
    endcase
  assign n11963_o = n11950_o[31:16];
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11954_o)
      3'b100: n11965_o = n11963_o;
      3'b010: n11965_o = 16'bX;
      3'b001: n11965_o = 16'bX;
      default: n11965_o = 16'bX;
    endcase
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11954_o)
      3'b100: n11966_o = n11951_o;
      3'b010: n11966_o = n11942_o;
      3'b001: n11966_o = n11936_o;
      default: n11966_o = n11928_o;
    endcase
  /* TG68K_ALU.vhd:809:38  */
  assign n11967_o = exe_opcode[8];
  /* TG68K_ALU.vhd:810:44  */
  assign n11968_o = alu[0];
  /* TG68K_ALU.vhd:809:25  */
  assign n11969_o = n11967_o ? n11968_o : n11966_o;
  /* TG68K_ALU.vhd:812:31  */
  assign n11971_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:813:40  */
  assign n11972_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:815:69  */
  assign n11973_o = result_bs[7:0];
  /* TG68K_ALU.vhd:815:94  */
  assign n11974_o = result_bs[16:9];
  /* TG68K_ALU.vhd:815:82  */
  assign n11975_o = n11973_o | n11974_o;
  /* TG68K_ALU.vhd:816:58  */
  assign n11976_o = result_bs[8];
  /* TG68K_ALU.vhd:816:74  */
  assign n11977_o = result_bs[17];
  /* TG68K_ALU.vhd:816:62  */
  assign n11978_o = n11976_o | n11977_o;
  /* TG68K_ALU.vhd:814:33  */
  assign n11980_o = n11972_o == 2'b00;
  /* TG68K_ALU.vhd:818:70  */
  assign n11981_o = result_bs[15:0];
  /* TG68K_ALU.vhd:818:96  */
  assign n11982_o = result_bs[32:17];
  /* TG68K_ALU.vhd:818:84  */
  assign n11983_o = n11981_o | n11982_o;
  /* TG68K_ALU.vhd:819:58  */
  assign n11984_o = result_bs[16];
  /* TG68K_ALU.vhd:819:75  */
  assign n11985_o = result_bs[33];
  /* TG68K_ALU.vhd:819:63  */
  assign n11986_o = n11984_o | n11985_o;
  /* TG68K_ALU.vhd:817:33  */
  assign n11988_o = n11972_o == 2'b01;
  /* TG68K_ALU.vhd:817:42  */
  assign n11990_o = n11972_o == 2'b11;
  /* TG68K_ALU.vhd:817:42  */
  assign n11991_o = n11988_o | n11990_o;
  /* TG68K_ALU.vhd:821:57  */
  assign n11992_o = result_bs[31:0];
  /* TG68K_ALU.vhd:821:83  */
  assign n11993_o = result_bs[64:33];
  /* TG68K_ALU.vhd:821:71  */
  assign n11994_o = n11992_o | n11993_o;
  /* TG68K_ALU.vhd:822:58  */
  assign n11995_o = result_bs[32];
  /* TG68K_ALU.vhd:822:75  */
  assign n11996_o = result_bs[65];
  /* TG68K_ALU.vhd:822:63  */
  assign n11997_o = n11995_o | n11996_o;
  /* TG68K_ALU.vhd:820:33  */
  assign n11999_o = n11972_o == 2'b10;
  assign n12000_o = {n11999_o, n11991_o, n11980_o};
  assign n12001_o = n11983_o[7:0];
  assign n12002_o = n11994_o[7:0];
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n12000_o)
      3'b100: n12004_o = n12002_o;
      3'b010: n12004_o = n12001_o;
      3'b001: n12004_o = n11975_o;
      default: n12004_o = 8'bX;
    endcase
  assign n12005_o = n11983_o[15:8];
  assign n12006_o = n11994_o[15:8];
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n12000_o)
      3'b100: n12008_o = n12006_o;
      3'b010: n12008_o = n12005_o;
      3'b001: n12008_o = 8'bX;
      default: n12008_o = 8'bX;
    endcase
  assign n12009_o = n11994_o[31:16];
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n12000_o)
      3'b100: n12011_o = n12009_o;
      3'b010: n12011_o = 16'bX;
      3'b001: n12011_o = 16'bX;
      default: n12011_o = 16'bX;
    endcase
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n12000_o)
      3'b100: n12012_o = n11997_o;
      3'b010: n12012_o = n11986_o;
      3'b001: n12012_o = n11978_o;
      default: n12012_o = n11928_o;
    endcase
  /* TG68K_ALU.vhd:826:38  */
  assign n12013_o = exe_opcode[8];
  /* TG68K_ALU.vhd:826:41  */
  assign n12014_o = ~n12013_o;
  /* TG68K_ALU.vhd:827:49  */
  assign n12015_o = result_bs[63:32];
  /* TG68K_ALU.vhd:829:49  */
  assign n12016_o = result_bs[31:0];
  /* TG68K_ALU.vhd:826:25  */
  assign n12017_o = n12014_o ? n12015_o : n12016_o;
  assign n12018_o = {n12011_o, n12008_o, n12004_o};
  /* TG68K_ALU.vhd:812:17  */
  assign n12019_o = n11971_o ? n12018_o : n12017_o;
  /* TG68K_ALU.vhd:812:17  */
  assign n12020_o = n11971_o ? n12012_o : n11928_o;
  assign n12021_o = {n11965_o, n11962_o, n11958_o};
  /* TG68K_ALU.vhd:795:17  */
  assign n12022_o = n11930_o ? n12021_o : n12019_o;
  /* TG68K_ALU.vhd:795:17  */
  assign n12024_o = n11930_o ? n11969_o : n12020_o;
  /* TG68K_ALU.vhd:795:17  */
  assign n12025_o = n11930_o ? n11931_o : bs_c;
  /* TG68K_ALU.vhd:833:29  */
  assign n12027_o = bs_shift == 6'b000000;
  /* TG68K_ALU.vhd:834:36  */
  assign n12029_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:835:46  */
  assign n12030_o = n12945_q[4];
  /* TG68K_ALU.vhd:834:25  */
  assign n12032_o = n12029_o ? n12030_o : 1'b0;
  /* TG68K_ALU.vhd:839:38  */
  assign n12033_o = n12945_q[4];
  /* TG68K_ALU.vhd:833:17  */
  assign n12035_o = n12027_o ? 1'b0 : n11908_o;
  /* TG68K_ALU.vhd:833:17  */
  assign n12036_o = n12027_o ? n12032_o : n12024_o;
  /* TG68K_ALU.vhd:833:17  */
  assign n12037_o = n12027_o ? n12033_o : n12025_o;
  /* TG68K_ALU.vhd:848:45  */
  assign n12039_o = bs_shift == 6'b111111;
  /* TG68K_ALU.vhd:850:48  */
  assign n12041_o = $unsigned(bs_shift) > $unsigned(6'b110101);
  /* TG68K_ALU.vhd:851:66  */
  assign n12043_o = bs_shift - 6'b110110;
  /* TG68K_ALU.vhd:852:48  */
  assign n12045_o = $unsigned(bs_shift) > $unsigned(6'b101100);
  /* TG68K_ALU.vhd:853:66  */
  assign n12047_o = bs_shift - 6'b101101;
  /* TG68K_ALU.vhd:854:48  */
  assign n12049_o = $unsigned(bs_shift) > $unsigned(6'b100011);
  /* TG68K_ALU.vhd:855:66  */
  assign n12051_o = bs_shift - 6'b100100;
  /* TG68K_ALU.vhd:856:48  */
  assign n12053_o = $unsigned(bs_shift) > $unsigned(6'b011010);
  /* TG68K_ALU.vhd:857:66  */
  assign n12055_o = bs_shift - 6'b011011;
  /* TG68K_ALU.vhd:858:48  */
  assign n12057_o = $unsigned(bs_shift) > $unsigned(6'b010001);
  /* TG68K_ALU.vhd:859:66  */
  assign n12059_o = bs_shift - 6'b010010;
  /* TG68K_ALU.vhd:860:48  */
  assign n12061_o = $unsigned(bs_shift) > $unsigned(6'b001000);
  /* TG68K_ALU.vhd:861:66  */
  assign n12063_o = bs_shift - 6'b001001;
  /* TG68K_ALU.vhd:860:33  */
  assign n12064_o = n12061_o ? n12063_o : bs_shift;
  /* TG68K_ALU.vhd:858:33  */
  assign n12065_o = n12057_o ? n12059_o : n12064_o;
  /* TG68K_ALU.vhd:856:33  */
  assign n12066_o = n12053_o ? n12055_o : n12065_o;
  /* TG68K_ALU.vhd:854:33  */
  assign n12067_o = n12049_o ? n12051_o : n12066_o;
  /* TG68K_ALU.vhd:852:33  */
  assign n12068_o = n12045_o ? n12047_o : n12067_o;
  /* TG68K_ALU.vhd:850:33  */
  assign n12069_o = n12041_o ? n12043_o : n12068_o;
  /* TG68K_ALU.vhd:848:33  */
  assign n12071_o = n12039_o ? 6'b000000 : n12069_o;
  /* TG68K_ALU.vhd:847:25  */
  assign n12073_o = ring == 6'b001001;
  /* TG68K_ALU.vhd:866:45  */
  assign n12075_o = $unsigned(bs_shift) > $unsigned(6'b110010);
  /* TG68K_ALU.vhd:867:66  */
  assign n12077_o = bs_shift - 6'b110011;
  /* TG68K_ALU.vhd:868:48  */
  assign n12079_o = $unsigned(bs_shift) > $unsigned(6'b100001);
  /* TG68K_ALU.vhd:869:66  */
  assign n12081_o = bs_shift - 6'b100010;
  /* TG68K_ALU.vhd:870:48  */
  assign n12083_o = $unsigned(bs_shift) > $unsigned(6'b010000);
  /* TG68K_ALU.vhd:871:66  */
  assign n12085_o = bs_shift - 6'b010001;
  /* TG68K_ALU.vhd:870:33  */
  assign n12086_o = n12083_o ? n12085_o : bs_shift;
  /* TG68K_ALU.vhd:868:33  */
  assign n12087_o = n12079_o ? n12081_o : n12086_o;
  /* TG68K_ALU.vhd:866:33  */
  assign n12088_o = n12075_o ? n12077_o : n12087_o;
  /* TG68K_ALU.vhd:865:25  */
  assign n12090_o = ring == 6'b010001;
  /* TG68K_ALU.vhd:876:45  */
  assign n12092_o = $unsigned(bs_shift) > $unsigned(6'b100000);
  /* TG68K_ALU.vhd:877:66  */
  assign n12094_o = bs_shift - 6'b100001;
  /* TG68K_ALU.vhd:876:33  */
  assign n12095_o = n12092_o ? n12094_o : bs_shift;
  /* TG68K_ALU.vhd:875:25  */
  assign n12097_o = ring == 6'b100001;
  /* TG68K_ALU.vhd:881:74  */
  assign n12098_o = bs_shift[2:0];
  /* TG68K_ALU.vhd:881:64  */
  assign n12100_o = {3'b000, n12098_o};
  /* TG68K_ALU.vhd:881:25  */
  assign n12102_o = ring == 6'b001000;
  /* TG68K_ALU.vhd:882:74  */
  assign n12103_o = bs_shift[3:0];
  /* TG68K_ALU.vhd:882:64  */
  assign n12105_o = {2'b00, n12103_o};
  /* TG68K_ALU.vhd:882:25  */
  assign n12107_o = ring == 6'b010000;
  /* TG68K_ALU.vhd:883:74  */
  assign n12108_o = bs_shift[4:0];
  /* TG68K_ALU.vhd:883:64  */
  assign n12110_o = {1'b0, n12108_o};
  /* TG68K_ALU.vhd:883:25  */
  assign n12112_o = ring == 6'b100000;
  assign n12113_o = {n12112_o, n12107_o, n12102_o, n12097_o, n12090_o, n12073_o};
  /* TG68K_ALU.vhd:846:17  */
  always @*
    case (n12113_o)
      6'b100000: n12115_o = n12110_o;
      6'b010000: n12115_o = n12105_o;
      6'b001000: n12115_o = n12100_o;
      6'b000100: n12115_o = n12095_o;
      6'b000010: n12115_o = n12088_o;
      6'b000001: n12115_o = n12071_o;
      default: n12115_o = 6'b000000;
    endcase
  /* TG68K_ALU.vhd:888:30  */
  assign n12116_o = exe_opcode[8];
  /* TG68K_ALU.vhd:888:33  */
  assign n12117_o = ~n12116_o;
  /* TG68K_ALU.vhd:889:39  */
  assign n12118_o = ring - bs_shift_mod;
  /* TG68K_ALU.vhd:888:17  */
  assign n12119_o = n12117_o ? n12118_o : bs_shift_mod;
  /* TG68K_ALU.vhd:891:28  */
  assign n12120_o = rot_bits[1];
  /* TG68K_ALU.vhd:891:31  */
  assign n12121_o = ~n12120_o;
  /* TG68K_ALU.vhd:892:38  */
  assign n12122_o = exe_opcode[8];
  /* TG68K_ALU.vhd:892:41  */
  assign n12123_o = ~n12122_o;
  /* TG68K_ALU.vhd:893:45  */
  assign n12125_o = 6'b100000 - bs_shift_mod;
  /* TG68K_ALU.vhd:892:25  */
  assign n12126_o = n12123_o ? n12125_o : n12119_o;
  /* TG68K_ALU.vhd:895:37  */
  assign n12127_o = bs_shift == ring;
  /* TG68K_ALU.vhd:896:46  */
  assign n12128_o = exe_opcode[8];
  /* TG68K_ALU.vhd:896:49  */
  assign n12129_o = ~n12128_o;
  /* TG68K_ALU.vhd:897:53  */
  assign n12131_o = 6'b100000 - ring;
  /* TG68K_ALU.vhd:896:33  */
  assign n12132_o = n12129_o ? n12131_o : ring;
  /* TG68K_ALU.vhd:895:25  */
  assign n12133_o = n12127_o ? n12132_o : n12126_o;
  /* TG68K_ALU.vhd:902:37  */
  assign n12134_o = $unsigned(bs_shift) > $unsigned(ring);
  /* TG68K_ALU.vhd:903:46  */
  assign n12135_o = exe_opcode[8];
  /* TG68K_ALU.vhd:903:49  */
  assign n12136_o = ~n12135_o;
  /* TG68K_ALU.vhd:907:55  */
  assign n12138_o = ring + 6'b000001;
  /* TG68K_ALU.vhd:903:33  */
  assign n12140_o = n12136_o ? 6'b000000 : n12138_o;
  /* TG68K_ALU.vhd:891:17  */
  assign n12142_o = n12146_o ? 1'b0 : n12036_o;
  /* TG68K_ALU.vhd:902:25  */
  assign n12143_o = n12134_o ? n12140_o : n12133_o;
  /* TG68K_ALU.vhd:902:25  */
  assign n12144_o = n12136_o & n12134_o;
  /* TG68K_ALU.vhd:891:17  */
  assign n12145_o = n12121_o ? n12143_o : n12119_o;
  /* TG68K_ALU.vhd:891:17  */
  assign n12146_o = n12144_o & n12121_o;
  /* TG68K_ALU.vhd:915:50  */
  assign n12147_o = asr_sign[31:0];
  /* TG68K_ALU.vhd:915:74  */
  assign n12148_o = hot_msb[31:0];
  /* TG68K_ALU.vhd:915:64  */
  assign n12149_o = n12147_o | n12148_o;
  assign n12151_o = n12150_o[0];
  /* TG68K_ALU.vhd:916:28  */
  assign n12153_o = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:916:48  */
  assign n12154_o = exe_opcode[8];
  /* TG68K_ALU.vhd:916:51  */
  assign n12155_o = ~n12154_o;
  /* TG68K_ALU.vhd:916:34  */
  assign n12156_o = n12155_o & n12153_o;
  /* TG68K_ALU.vhd:916:56  */
  assign n12157_o = msb & n12156_o;
  /* TG68K_ALU.vhd:917:49  */
  assign n12158_o = asr_sign[32:1];
  /* TG68K_ALU.vhd:917:38  */
  assign n12159_o = alu | n12158_o;
  /* TG68K_ALU.vhd:918:37  */
  assign n12160_o = $unsigned(bs_shift) > $unsigned(ring);
  /* TG68K_ALU.vhd:916:17  */
  assign n12162_o = n12164_o ? 1'b1 : n12142_o;
  /* TG68K_ALU.vhd:916:17  */
  assign n12164_o = n12160_o & n12157_o;
  /* TG68K_ALU.vhd:923:43  */
  assign n12166_o = {1'b0, op1out};
  /* TG68K_ALU.vhd:924:32  */
  assign n12167_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:926:46  */
  assign n12168_o = op1out[7];
  /* TG68K_ALU.vhd:929:44  */
  assign n12172_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:930:59  */
  assign n12173_o = n12945_q[4];
  assign n12174_o = n12169_o[0];
  /* TG68K_ALU.vhd:929:33  */
  assign n12175_o = n12172_o ? n12173_o : n12174_o;
  assign n12176_o = n12169_o[23:1];
  /* TG68K_ALU.vhd:925:25  */
  assign n12178_o = n12167_o == 2'b00;
  /* TG68K_ALU.vhd:933:46  */
  assign n12179_o = op1out[15];
  /* TG68K_ALU.vhd:936:44  */
  assign n12183_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:937:60  */
  assign n12184_o = n12945_q[4];
  assign n12185_o = n12180_o[0];
  /* TG68K_ALU.vhd:936:33  */
  assign n12186_o = n12183_o ? n12184_o : n12185_o;
  assign n12187_o = n12180_o[15:1];
  /* TG68K_ALU.vhd:932:25  */
  assign n12189_o = n12167_o == 2'b01;
  /* TG68K_ALU.vhd:932:34  */
  assign n12191_o = n12167_o == 2'b11;
  /* TG68K_ALU.vhd:932:34  */
  assign n12192_o = n12189_o | n12191_o;
  /* TG68K_ALU.vhd:940:46  */
  assign n12193_o = op1out[31];
  /* TG68K_ALU.vhd:941:44  */
  assign n12195_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:942:60  */
  assign n12196_o = n12945_q[4];
  assign n12197_o = n12166_o[32];
  /* TG68K_ALU.vhd:941:33  */
  assign n12198_o = n12195_o ? n12196_o : n12197_o;
  /* TG68K_ALU.vhd:939:25  */
  assign n12200_o = n12167_o == 2'b10;
  assign n12201_o = {n12200_o, n12192_o, n12178_o};
  assign n12202_o = n12166_o[8];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12203_o = n12202_o;
      3'b010: n12203_o = n12202_o;
      3'b001: n12203_o = n12175_o;
      default: n12203_o = n12202_o;
    endcase
  assign n12204_o = n12176_o[6:0];
  assign n12205_o = n12166_o[15:9];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12206_o = n12205_o;
      3'b010: n12206_o = n12205_o;
      3'b001: n12206_o = n12204_o;
      default: n12206_o = n12205_o;
    endcase
  assign n12207_o = n12176_o[7];
  assign n12208_o = n12166_o[16];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12209_o = n12208_o;
      3'b010: n12209_o = n12186_o;
      3'b001: n12209_o = n12207_o;
      default: n12209_o = n12208_o;
    endcase
  assign n12210_o = n12176_o[22:8];
  assign n12211_o = n12166_o[31:17];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12212_o = n12211_o;
      3'b010: n12212_o = n12187_o;
      3'b001: n12212_o = n12210_o;
      default: n12212_o = n12211_o;
    endcase
  assign n12213_o = n12166_o[32];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12214_o = n12198_o;
      3'b010: n12214_o = n12213_o;
      3'b001: n12214_o = n12213_o;
      default: n12214_o = n12213_o;
    endcase
  assign n12216_o = n12166_o[7:0];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12220_o = n12193_o;
      3'b010: n12220_o = n12179_o;
      3'b001: n12220_o = n12168_o;
      default: n12220_o = msb;
    endcase
  assign n12221_o = n12170_o[7:0];
  assign n12222_o = n12159_o[15:8];
  assign n12223_o = alu[15:8];
  /* TG68K_ALU.vhd:916:17  */
  assign n12224_o = n12157_o ? n12222_o : n12223_o;
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12225_o = n12224_o;
      3'b010: n12225_o = n12224_o;
      3'b001: n12225_o = n12221_o;
      default: n12225_o = n12224_o;
    endcase
  assign n12226_o = n12170_o[23:8];
  assign n12227_o = n12159_o[31:16];
  assign n12228_o = alu[31:16];
  /* TG68K_ALU.vhd:916:17  */
  assign n12229_o = n12157_o ? n12227_o : n12228_o;
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12201_o)
      3'b100: n12230_o = n12229_o;
      3'b010: n12230_o = 16'b0000000000000000;
      3'b001: n12230_o = n12226_o;
      default: n12230_o = n12229_o;
    endcase
  assign n12234_o = n12159_o[7:0];
  assign n12235_o = alu[7:0];
  /* TG68K_ALU.vhd:916:17  */
  assign n12236_o = n12157_o ? n12234_o : n12235_o;
  /* TG68K_ALU.vhd:946:71  */
  assign n12238_o = {33'b000000000000000000000000000000000, vector};
  /* TG68K_ALU.vhd:946:84  */
  assign n12239_o = {25'b0, bit_nr};  //  uext
  /* TG68K_ALU.vhd:946:80  */
  assign n12240_o = {1'b0, n12239_o};  //  uext
  /* TG68K_ALU.vhd:946:80  */
  assign n12241_o = n12238_o << n12240_o;
  /* TG68K_ALU.vhd:957:24  */
  assign n12245_o = exec[17];
  /* TG68K_ALU.vhd:958:58  */
  assign n12246_o = last_data_read[7:0];
  /* TG68K_ALU.vhd:958:40  */
  assign n12247_o = n12945_q & n12246_o;
  /* TG68K_ALU.vhd:959:27  */
  assign n12248_o = exec[18];
  /* TG68K_ALU.vhd:960:58  */
  assign n12249_o = last_data_read[7:0];
  /* TG68K_ALU.vhd:960:40  */
  assign n12250_o = n12945_q ^ n12249_o;
  /* TG68K_ALU.vhd:961:27  */
  assign n12251_o = exec[19];
  /* TG68K_ALU.vhd:962:57  */
  assign n12252_o = last_data_read[7:0];
  /* TG68K_ALU.vhd:962:40  */
  assign n12253_o = n12945_q | n12252_o;
  /* TG68K_ALU.vhd:964:40  */
  assign n12254_o = op2out[7:0];
  /* TG68K_ALU.vhd:961:17  */
  assign n12255_o = n12251_o ? n12253_o : n12254_o;
  /* TG68K_ALU.vhd:959:17  */
  assign n12256_o = n12248_o ? n12250_o : n12255_o;
  /* TG68K_ALU.vhd:957:17  */
  assign n12257_o = n12245_o ? n12247_o : n12256_o;
  /* TG68K_ALU.vhd:971:24  */
  assign n12258_o = exec[28];
  /* TG68K_ALU.vhd:971:50  */
  assign n12259_o = n12945_q[2];
  /* TG68K_ALU.vhd:971:53  */
  assign n12260_o = ~n12259_o;
  /* TG68K_ALU.vhd:971:41  */
  assign n12261_o = n12260_o & n12258_o;
  /* TG68K_ALU.vhd:973:28  */
  assign n12262_o = op1in[7:0];
  /* TG68K_ALU.vhd:973:40  */
  assign n12264_o = n12262_o == 8'b00000000;
  /* TG68K_ALU.vhd:975:33  */
  assign n12266_o = op1in[15:8];
  /* TG68K_ALU.vhd:975:46  */
  assign n12268_o = n12266_o == 8'b00000000;
  /* TG68K_ALU.vhd:977:41  */
  assign n12270_o = op1in[31:16];
  /* TG68K_ALU.vhd:977:55  */
  assign n12272_o = n12270_o == 16'b0000000000000000;
  /* TG68K_ALU.vhd:977:33  */
  assign n12275_o = n12272_o ? 1'b1 : 1'b0;
  assign n12276_o = {n12275_o, 1'b1};
  /* TG68K_ALU.vhd:975:25  */
  assign n12278_o = n12268_o ? n12276_o : 2'b00;
  assign n12279_o = {n12278_o, 1'b1};
  /* TG68K_ALU.vhd:973:17  */
  assign n12281_o = n12264_o ? n12279_o : 3'b000;
  /* TG68K_ALU.vhd:971:17  */
  assign n12283_o = n12261_o ? 3'b000 : n12281_o;
  /* TG68K_ALU.vhd:984:32  */
  assign n12286_o = exe_datatype == 2'b00;
  /* TG68K_ALU.vhd:985:43  */
  assign n12287_o = op1in[7];
  /* TG68K_ALU.vhd:985:53  */
  assign n12288_o = flag_z[0];
  /* TG68K_ALU.vhd:985:46  */
  assign n12289_o = {n12287_o, n12288_o};
  /* TG68K_ALU.vhd:985:67  */
  assign n12290_o = addsub_ofl[0];
  /* TG68K_ALU.vhd:985:56  */
  assign n12291_o = {n12289_o, n12290_o};
  /* TG68K_ALU.vhd:985:76  */
  assign n12292_o = n10188_o[0];
  /* TG68K_ALU.vhd:985:70  */
  assign n12293_o = {n12291_o, n12292_o};
  /* TG68K_ALU.vhd:986:32  */
  assign n12294_o = exec[12];
  /* TG68K_ALU.vhd:986:53  */
  assign n12295_o = exec[13];
  /* TG68K_ALU.vhd:986:46  */
  assign n12296_o = n12294_o | n12295_o;
  assign n12297_o = {vflag_a, bcd_a_carry};
  assign n12298_o = n12293_o[1:0];
  /* TG68K_ALU.vhd:986:25  */
  assign n12299_o = n12296_o ? n12297_o : n12298_o;
  assign n12300_o = n12293_o[3:2];
  /* TG68K_ALU.vhd:990:35  */
  assign n12302_o = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:990:48  */
  assign n12303_o = exec[10];
  /* TG68K_ALU.vhd:990:41  */
  assign n12304_o = n12302_o | n12303_o;
  /* TG68K_ALU.vhd:991:43  */
  assign n12305_o = op1in[31];
  /* TG68K_ALU.vhd:991:54  */
  assign n12306_o = flag_z[2];
  /* TG68K_ALU.vhd:991:47  */
  assign n12307_o = {n12305_o, n12306_o};
  /* TG68K_ALU.vhd:991:68  */
  assign n12308_o = addsub_ofl[2];
  /* TG68K_ALU.vhd:991:57  */
  assign n12309_o = {n12307_o, n12308_o};
  /* TG68K_ALU.vhd:991:77  */
  assign n12310_o = n10188_o[2];
  /* TG68K_ALU.vhd:991:71  */
  assign n12311_o = {n12309_o, n12310_o};
  /* TG68K_ALU.vhd:993:43  */
  assign n12312_o = op1in[15];
  /* TG68K_ALU.vhd:993:54  */
  assign n12313_o = flag_z[1];
  /* TG68K_ALU.vhd:993:47  */
  assign n12314_o = {n12312_o, n12313_o};
  /* TG68K_ALU.vhd:993:68  */
  assign n12315_o = addsub_ofl[1];
  /* TG68K_ALU.vhd:993:57  */
  assign n12316_o = {n12314_o, n12315_o};
  /* TG68K_ALU.vhd:993:77  */
  assign n12317_o = n10188_o[1];
  /* TG68K_ALU.vhd:993:71  */
  assign n12318_o = {n12316_o, n12317_o};
  /* TG68K_ALU.vhd:990:17  */
  assign n12319_o = n12304_o ? n12311_o : n12318_o;
  assign n12320_o = {n12300_o, n12299_o};
  /* TG68K_ALU.vhd:984:17  */
  assign n12321_o = n12286_o ? n12320_o : n12319_o;
  /* TG68K_ALU.vhd:1000:40  */
  assign n12323_o = exec[59];
  /* TG68K_ALU.vhd:1000:55  */
  assign n12324_o = n12323_o | set_stop;
  /* TG68K_ALU.vhd:1003:40  */
  assign n12327_o = exec[60];
  /* TG68K_ALU.vhd:1007:40  */
  assign n12330_o = exec[9];
  /* TG68K_ALU.vhd:1007:66  */
  assign n12331_o = ~decodeopc;
  /* TG68K_ALU.vhd:1007:53  */
  assign n12332_o = n12331_o & n12330_o;
  /* TG68K_ALU.vhd:1008:65  */
  assign n12333_o = set_flags[3];
  /* TG68K_ALU.vhd:1008:69  */
  assign n12334_o = n12333_o ^ rot_rot;
  /* TG68K_ALU.vhd:1008:82  */
  assign n12335_o = n12334_o | asl_vflag;
  /* TG68K_ALU.vhd:1007:33  */
  assign n12337_o = n12332_o ? n12335_o : 1'b0;
  /* TG68K_ALU.vhd:1012:40  */
  assign n12338_o = exec[51];
  /* TG68K_ALU.vhd:1015:56  */
  assign n12340_o = micro_state == 7'b0110011;
  /* TG68K_ALU.vhd:1017:62  */
  assign n12341_o = exe_opcode[8];
  /* TG68K_ALU.vhd:1017:65  */
  assign n12342_o = ~n12341_o;
  /* TG68K_ALU.vhd:1019:92  */
  assign n12343_o = reg_qa[31];
  /* TG68K_ALU.vhd:1019:82  */
  assign n12344_o = ~n12343_o;
  /* TG68K_ALU.vhd:1019:81  */
  assign n12346_o = {1'b0, n12344_o};
  /* TG68K_ALU.vhd:1019:96  */
  assign n12348_o = {n12346_o, 2'b00};
  /* TG68K_ALU.vhd:1017:49  */
  assign n12350_o = n12342_o ? n12348_o : 4'b0100;
  assign n12351_o = data_read[3:0];
  assign n12352_o = data_read[3:0];
  assign n12353_o = n12945_q[3:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12354_o = n12324_o ? n12352_o : n12353_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12355_o = n12327_o ? n12351_o : n12354_o;
  /* TG68K_ALU.vhd:1015:41  */
  assign n12356_o = n12340_o ? n12350_o : n12355_o;
  /* TG68K_ALU.vhd:1024:43  */
  assign n12357_o = exec[49];
  /* TG68K_ALU.vhd:1024:53  */
  assign n12358_o = ~n12357_o;
  /* TG68K_ALU.vhd:1025:61  */
  assign n12359_o = n12945_q[3:0];
  /* TG68K_ALU.vhd:1026:48  */
  assign n12360_o = exec[3];
  /* TG68K_ALU.vhd:1027:70  */
  assign n12361_o = set_flags[0];
  /* TG68K_ALU.vhd:1028:51  */
  assign n12362_o = exec[9];
  /* TG68K_ALU.vhd:1028:76  */
  assign n12364_o = rot_bits != 2'b11;
  /* TG68K_ALU.vhd:1028:64  */
  assign n12365_o = n12364_o & n12362_o;
  /* TG68K_ALU.vhd:1028:91  */
  assign n12366_o = exec[23];
  /* TG68K_ALU.vhd:1028:100  */
  assign n12367_o = ~n12366_o;
  /* TG68K_ALU.vhd:1028:83  */
  assign n12368_o = n12367_o & n12365_o;
  /* TG68K_ALU.vhd:1030:51  */
  assign n12369_o = exec[81];
  assign n12370_o = data_read[4];
  assign n12371_o = data_read[4];
  assign n12372_o = n12945_q[4];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12373_o = n12324_o ? n12371_o : n12372_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12374_o = n12327_o ? n12370_o : n12373_o;
  /* TG68K_ALU.vhd:1030:41  */
  assign n12375_o = n12369_o ? bs_x : n12374_o;
  /* TG68K_ALU.vhd:1028:41  */
  assign n12376_o = n12368_o ? rot_x : n12375_o;
  /* TG68K_ALU.vhd:1026:41  */
  assign n12377_o = n12360_o ? n12361_o : n12376_o;
  /* TG68K_ALU.vhd:1034:49  */
  assign n12378_o = exec[8];
  /* TG68K_ALU.vhd:1034:65  */
  assign n12379_o = exec[86];
  /* TG68K_ALU.vhd:1034:58  */
  assign n12380_o = n12378_o | n12379_o;
  /* TG68K_ALU.vhd:1036:51  */
  assign n12381_o = exec[21];
  /* TG68K_ALU.vhd:1036:65  */
  assign n12383_o = 1'b1 & n12381_o;
  /* TG68K_ALU.vhd:1039:65  */
  assign n12385_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1039:74  */
  assign n12387_o = n12385_o | 1'b0;
  /* TG68K_ALU.vhd:1040:83  */
  assign n12388_o = op1in[15];
  /* TG68K_ALU.vhd:1040:94  */
  assign n12389_o = flag_z[1];
  /* TG68K_ALU.vhd:1040:87  */
  assign n12390_o = {n12388_o, n12389_o};
  /* TG68K_ALU.vhd:1040:97  */
  assign n12392_o = {n12390_o, 2'b00};
  /* TG68K_ALU.vhd:1042:83  */
  assign n12393_o = op1in[31];
  /* TG68K_ALU.vhd:1042:94  */
  assign n12394_o = flag_z[2];
  /* TG68K_ALU.vhd:1042:87  */
  assign n12395_o = {n12393_o, n12394_o};
  /* TG68K_ALU.vhd:1042:97  */
  assign n12397_o = {n12395_o, 2'b00};
  /* TG68K_ALU.vhd:1039:49  */
  assign n12398_o = n12387_o ? n12392_o : n12397_o;
  /* TG68K_ALU.vhd:1037:49  */
  assign n12399_o = v_flag ? 4'b1010 : n12398_o;
  /* TG68K_ALU.vhd:1044:51  */
  assign n12400_o = exec[68];
  /* TG68K_ALU.vhd:1044:72  */
  assign n12402_o = 1'b1 & n12400_o;
  /* TG68K_ALU.vhd:1045:70  */
  assign n12403_o = set_flags[3];
  /* TG68K_ALU.vhd:1046:70  */
  assign n12404_o = set_flags[2];
  /* TG68K_ALU.vhd:1046:83  */
  assign n12405_o = n12945_q[2];
  /* TG68K_ALU.vhd:1046:74  */
  assign n12406_o = n12404_o & n12405_o;
  /* TG68K_ALU.vhd:1049:51  */
  assign n12409_o = exec[67];
  /* TG68K_ALU.vhd:1049:71  */
  assign n12411_o = 1'b1 & n12409_o;
  /* TG68K_ALU.vhd:1050:70  */
  assign n12412_o = set_flags[3];
  /* TG68K_ALU.vhd:1051:70  */
  assign n12413_o = set_flags[2];
  /* TG68K_ALU.vhd:1054:51  */
  assign n12415_o = exec[5];
  /* TG68K_ALU.vhd:1054:70  */
  assign n12416_o = exec[6];
  /* TG68K_ALU.vhd:1054:63  */
  assign n12417_o = n12415_o | n12416_o;
  /* TG68K_ALU.vhd:1054:90  */
  assign n12418_o = exec[7];
  /* TG68K_ALU.vhd:1054:83  */
  assign n12419_o = n12417_o | n12418_o;
  /* TG68K_ALU.vhd:1054:110  */
  assign n12420_o = exec[0];
  /* TG68K_ALU.vhd:1054:103  */
  assign n12421_o = n12419_o | n12420_o;
  /* TG68K_ALU.vhd:1054:131  */
  assign n12422_o = exec[1];
  /* TG68K_ALU.vhd:1054:124  */
  assign n12423_o = n12421_o | n12422_o;
  /* TG68K_ALU.vhd:1054:153  */
  assign n12424_o = exec[15];
  /* TG68K_ALU.vhd:1054:146  */
  assign n12425_o = n12423_o | n12424_o;
  /* TG68K_ALU.vhd:1054:174  */
  assign n12426_o = exec[75];
  /* TG68K_ALU.vhd:1054:167  */
  assign n12427_o = n12425_o | n12426_o;
  /* TG68K_ALU.vhd:1054:194  */
  assign n12428_o = exec[20];
  /* TG68K_ALU.vhd:1054:208  */
  assign n12430_o = 1'b1 & n12428_o;
  /* TG68K_ALU.vhd:1054:186  */
  assign n12431_o = n12427_o | n12430_o;
  /* TG68K_ALU.vhd:1057:56  */
  assign n12434_o = exec[75];
  assign n12435_o = set_flags[3];
  /* TG68K_ALU.vhd:1057:49  */
  assign n12436_o = n12434_o ? bf_nflag : n12435_o;
  assign n12437_o = set_flags[2];
  /* TG68K_ALU.vhd:1060:51  */
  assign n12438_o = exec[9];
  /* TG68K_ALU.vhd:1061:79  */
  assign n12439_o = set_flags[3:2];
  /* TG68K_ALU.vhd:1063:60  */
  assign n12441_o = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:1063:81  */
  assign n12442_o = set_flags[3];
  /* TG68K_ALU.vhd:1063:85  */
  assign n12443_o = n12442_o ^ rot_rot;
  /* TG68K_ALU.vhd:1063:98  */
  assign n12444_o = n12443_o | asl_vflag;
  /* TG68K_ALU.vhd:1063:66  */
  assign n12445_o = n12444_o & n12441_o;
  /* TG68K_ALU.vhd:1063:49  */
  assign n12448_o = n12445_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1068:51  */
  assign n12449_o = exec[81];
  /* TG68K_ALU.vhd:1069:79  */
  assign n12450_o = set_flags[3:2];
  /* TG68K_ALU.vhd:1072:51  */
  assign n12451_o = exec[14];
  /* TG68K_ALU.vhd:1073:61  */
  assign n12452_o = ~one_bit_in;
  /* TG68K_ALU.vhd:1074:51  */
  assign n12453_o = exec[87];
  /* TG68K_ALU.vhd:1079:63  */
  assign n12454_o = last_flags1[0];
  /* TG68K_ALU.vhd:1079:66  */
  assign n12455_o = ~n12454_o;
  /* TG68K_ALU.vhd:1080:74  */
  assign n12456_o = n12945_q[0];
  /* TG68K_ALU.vhd:1080:95  */
  assign n12457_o = set_flags[0];
  /* TG68K_ALU.vhd:1080:82  */
  assign n12458_o = ~n12457_o;
  /* TG68K_ALU.vhd:1080:116  */
  assign n12459_o = set_flags[2];
  /* TG68K_ALU.vhd:1080:103  */
  assign n12460_o = ~n12459_o;
  /* TG68K_ALU.vhd:1080:99  */
  assign n12461_o = n12458_o & n12460_o;
  /* TG68K_ALU.vhd:1080:78  */
  assign n12462_o = n12456_o | n12461_o;
  /* TG68K_ALU.vhd:1082:75  */
  assign n12463_o = n12945_q[0];
  /* TG68K_ALU.vhd:1082:92  */
  assign n12464_o = set_flags[0];
  /* TG68K_ALU.vhd:1082:79  */
  assign n12465_o = n12463_o ^ n12464_o;
  /* TG68K_ALU.vhd:1082:111  */
  assign n12466_o = n12945_q[2];
  /* TG68K_ALU.vhd:1082:102  */
  assign n12467_o = ~n12466_o;
  /* TG68K_ALU.vhd:1082:97  */
  assign n12468_o = n12465_o & n12467_o;
  /* TG68K_ALU.vhd:1082:132  */
  assign n12469_o = set_flags[2];
  /* TG68K_ALU.vhd:1082:119  */
  assign n12470_o = ~n12469_o;
  /* TG68K_ALU.vhd:1082:115  */
  assign n12471_o = n12468_o & n12470_o;
  /* TG68K_ALU.vhd:1079:49  */
  assign n12472_o = n12455_o ? n12462_o : n12471_o;
  /* TG68K_ALU.vhd:1085:66  */
  assign n12474_o = n12945_q[2];
  /* TG68K_ALU.vhd:1085:82  */
  assign n12475_o = set_flags[2];
  /* TG68K_ALU.vhd:1085:70  */
  assign n12476_o = n12474_o | n12475_o;
  /* TG68K_ALU.vhd:1086:76  */
  assign n12477_o = last_flags1[0];
  /* TG68K_ALU.vhd:1086:61  */
  assign n12478_o = ~n12477_o;
  /* TG68K_ALU.vhd:1087:51  */
  assign n12479_o = exec[31];
  /* TG68K_ALU.vhd:1088:64  */
  assign n12481_o = exe_datatype == 2'b01;
  /* TG68K_ALU.vhd:1089:75  */
  assign n12482_o = op1out[15];
  /* TG68K_ALU.vhd:1091:75  */
  assign n12483_o = op1out[31];
  /* TG68K_ALU.vhd:1088:49  */
  assign n12484_o = n12481_o ? n12482_o : n12483_o;
  /* TG68K_ALU.vhd:1093:58  */
  assign n12485_o = op1out[15:0];
  /* TG68K_ALU.vhd:1093:71  */
  assign n12487_o = n12485_o == 16'b0000000000000000;
  /* TG68K_ALU.vhd:1093:97  */
  assign n12489_o = exe_datatype == 2'b01;
  /* TG68K_ALU.vhd:1093:112  */
  assign n12490_o = op1out[31:16];
  /* TG68K_ALU.vhd:1093:126  */
  assign n12492_o = n12490_o == 16'b0000000000000000;
  /* TG68K_ALU.vhd:1093:103  */
  assign n12493_o = n12489_o | n12492_o;
  /* TG68K_ALU.vhd:1093:80  */
  assign n12494_o = n12493_o & n12487_o;
  /* TG68K_ALU.vhd:1093:49  */
  assign n12497_o = n12494_o ? 1'b1 : 1'b0;
  assign n12500_o = {n12484_o, n12497_o, 1'b0, 1'b0};
  assign n12501_o = data_read[3:0];
  assign n12502_o = data_read[3:0];
  assign n12503_o = n12945_q[3:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12504_o = n12324_o ? n12502_o : n12503_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12505_o = n12327_o ? n12501_o : n12504_o;
  /* TG68K_ALU.vhd:1087:41  */
  assign n12506_o = n12479_o ? n12500_o : n12505_o;
  assign n12507_o = {n12478_o, n12476_o, 1'b0, n12472_o};
  /* TG68K_ALU.vhd:1074:41  */
  assign n12508_o = n12453_o ? n12507_o : n12506_o;
  assign n12509_o = n12508_o[1:0];
  assign n12510_o = data_read[1:0];
  assign n12511_o = data_read[1:0];
  assign n12512_o = n12945_q[1:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12513_o = n12324_o ? n12511_o : n12512_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12514_o = n12327_o ? n12510_o : n12513_o;
  /* TG68K_ALU.vhd:1072:41  */
  assign n12515_o = n12451_o ? n12514_o : n12509_o;
  assign n12516_o = n12508_o[2];
  /* TG68K_ALU.vhd:1072:41  */
  assign n12517_o = n12451_o ? n12452_o : n12516_o;
  assign n12518_o = n12508_o[3];
  assign n12519_o = data_read[3];
  assign n12520_o = data_read[3];
  assign n12521_o = n12945_q[3];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12522_o = n12324_o ? n12520_o : n12521_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12523_o = n12327_o ? n12519_o : n12522_o;
  /* TG68K_ALU.vhd:1072:41  */
  assign n12524_o = n12451_o ? n12523_o : n12518_o;
  assign n12525_o = {n12524_o, n12517_o, n12515_o};
  assign n12526_o = {n12450_o, bs_v, bs_c};
  /* TG68K_ALU.vhd:1068:41  */
  assign n12527_o = n12449_o ? n12526_o : n12525_o;
  assign n12528_o = {n12439_o, n12448_o, rot_c};
  /* TG68K_ALU.vhd:1060:41  */
  assign n12529_o = n12438_o ? n12528_o : n12527_o;
  assign n12530_o = {n12436_o, n12437_o, 2'b00};
  /* TG68K_ALU.vhd:1054:41  */
  assign n12531_o = n12431_o ? n12530_o : n12529_o;
  assign n12532_o = {n12412_o, n12413_o, set_mv_flag, 1'b0};
  /* TG68K_ALU.vhd:1049:41  */
  assign n12533_o = n12411_o ? n12532_o : n12531_o;
  assign n12534_o = {n12403_o, n12406_o, 1'b0, 1'b0};
  /* TG68K_ALU.vhd:1044:41  */
  assign n12535_o = n12402_o ? n12534_o : n12533_o;
  /* TG68K_ALU.vhd:1036:41  */
  assign n12536_o = n12383_o ? n12399_o : n12535_o;
  /* TG68K_ALU.vhd:1034:41  */
  assign n12537_o = n12380_o ? set_flags : n12536_o;
  assign n12538_o = {n12377_o, n12537_o};
  assign n12539_o = data_read[4:0];
  assign n12540_o = data_read[4:0];
  assign n12541_o = n12945_q[4:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12542_o = n12324_o ? n12540_o : n12541_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12543_o = n12327_o ? n12539_o : n12542_o;
  /* TG68K_ALU.vhd:1024:33  */
  assign n12544_o = n12358_o ? n12538_o : n12543_o;
  /* TG68K_ALU.vhd:1024:33  */
  assign n12545_o = n12358_o ? n12359_o : last_flags1;
  assign n12546_o = n12544_o[3:0];
  /* TG68K_ALU.vhd:1014:33  */
  assign n12547_o = z_error ? n12356_o : n12546_o;
  assign n12548_o = n12544_o[4];
  assign n12549_o = data_read[4];
  assign n12550_o = data_read[4];
  assign n12551_o = n12945_q[4];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12552_o = n12324_o ? n12550_o : n12551_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12553_o = n12327_o ? n12549_o : n12552_o;
  /* TG68K_ALU.vhd:1014:33  */
  assign n12554_o = z_error ? n12553_o : n12548_o;
  /* TG68K_ALU.vhd:1014:33  */
  assign n12555_o = z_error ? last_flags1 : n12545_o;
  assign n12556_o = {n12554_o, n12547_o};
  assign n12557_o = ccrin[4:0];
  /* TG68K_ALU.vhd:1012:33  */
  assign n12558_o = n12338_o ? n12557_o : n12556_o;
  assign n12559_o = ccrin[7:5];
  assign n12560_o = data_read[7:5];
  assign n12561_o = data_read[7:5];
  assign n12562_o = n12945_q[7:5];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12563_o = n12324_o ? n12561_o : n12562_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12564_o = n12327_o ? n12560_o : n12563_o;
  /* TG68K_ALU.vhd:1012:33  */
  assign n12565_o = n12338_o ? n12559_o : n12564_o;
  /* TG68K_ALU.vhd:1012:33  */
  assign n12571_o = n12338_o ? last_flags1 : n12555_o;
  assign n12572_o = {n12565_o, n12558_o};
  /* TG68K_ALU.vhd:999:25  */
  assign n12574_o = clkena_lw ? n12571_o : last_flags1;
  /* TG68K_ALU.vhd:999:25  */
  assign n12575_o = clkena_lw ? n12337_o : asl_vflag;
  /* TG68K_ALU.vhd:997:25  */
  assign n12578_o = reset ? last_flags1 : n12574_o;
  /* TG68K_ALU.vhd:997:25  */
  assign n12579_o = reset ? asl_vflag : n12575_o;
  assign n12581_o = n12576_o[4:0];
  assign n12582_o = n12572_o[4:0];
  assign n12583_o = n12945_q[4:0];
  /* TG68K_ALU.vhd:999:25  */
  assign n12584_o = clkena_lw ? n12582_o : n12583_o;
  /* TG68K_ALU.vhd:997:25  */
  assign n12585_o = reset ? n12581_o : n12584_o;
  assign n12586_o = {3'b000, n12585_o};
  /* TG68K_ALU.vhd:1128:38  */
  assign n12593_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1129:59  */
  assign n12594_o = reg_qa[15];
  /* TG68K_ALU.vhd:1129:49  */
  assign n12595_o = n12594_o & signedop;
  /* TG68K_ALU.vhd:1129:33  */
  assign n12598_o = n12595_o ? 32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
  /* TG68K_ALU.vhd:1134:59  */
  assign n12599_o = op2out[15];
  /* TG68K_ALU.vhd:1134:49  */
  assign n12600_o = n12599_o & signedop;
  /* TG68K_ALU.vhd:1134:33  */
  assign n12603_o = n12600_o ? 32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
  /* TG68K_ALU.vhd:1140:63  */
  assign n12604_o = reg_qa[31:16];
  /* TG68K_ALU.vhd:1141:63  */
  assign n12605_o = op2out[31:16];
  /* TG68K_ALU.vhd:1142:59  */
  assign n12606_o = reg_qa[31];
  /* TG68K_ALU.vhd:1142:49  */
  assign n12607_o = n12606_o & signedop;
  /* TG68K_ALU.vhd:1142:33  */
  assign n12610_o = n12607_o ? 16'b1111111111111111 : 16'b0000000000000000;
  /* TG68K_ALU.vhd:1147:59  */
  assign n12611_o = op2out[31];
  /* TG68K_ALU.vhd:1147:49  */
  assign n12612_o = n12611_o & signedop;
  /* TG68K_ALU.vhd:1147:33  */
  assign n12615_o = n12612_o ? 16'b1111111111111111 : 16'b0000000000000000;
  assign n12616_o = {n12610_o, n12604_o};
  /* TG68K_ALU.vhd:1128:25  */
  assign n12617_o = n12593_o ? n12598_o : n12616_o;
  assign n12618_o = {n12615_o, n12605_o};
  /* TG68K_ALU.vhd:1128:25  */
  assign n12619_o = n12593_o ? n12603_o : n12618_o;
  /* TG68K_ALU.vhd:1153:62  */
  assign n12620_o = faktora[31:16];
  /* TG68K_ALU.vhd:1153:77  */
  assign n12621_o = {n12620_o, faktora};
  /* TG68K_ALU.vhd:1153:108  */
  assign n12622_o = reg_qa[15:0];
  /* TG68K_ALU.vhd:1153:100  */
  assign n12623_o = {n12621_o, n12622_o};
  /* TG68K_ALU.vhd:1153:133  */
  assign n12624_o = faktorb[31:16];
  /* TG68K_ALU.vhd:1153:148  */
  assign n12625_o = {n12624_o, faktorb};
  /* TG68K_ALU.vhd:1153:179  */
  assign n12626_o = op2out[15:0];
  /* TG68K_ALU.vhd:1153:171  */
  assign n12627_o = {n12625_o, n12626_o};
  /* TG68K_ALU.vhd:1153:123  */
  assign n12628_o = {64'b0, n12623_o};  //  uext
  /* TG68K_ALU.vhd:1153:123  */
  assign n12629_o = {64'b0, n12627_o};  //  uext
  /* TG68K_ALU.vhd:1153:123  */
  assign n12630_o = n12628_o * n12629_o; // umul
  /* TG68K_ALU.vhd:1201:32  */
  assign n12631_o = result_mulu[63:32];
  /* TG68K_ALU.vhd:1201:46  */
  assign n12633_o = n12631_o == 32'b00000000000000000000000000000000;
  /* TG68K_ALU.vhd:1201:72  */
  assign n12634_o = ~signedop;
  /* TG68K_ALU.vhd:1201:91  */
  assign n12635_o = result_mulu[31];
  /* TG68K_ALU.vhd:1201:95  */
  assign n12636_o = ~n12635_o;
  /* TG68K_ALU.vhd:1201:77  */
  assign n12637_o = n12634_o | n12636_o;
  /* TG68K_ALU.vhd:1201:59  */
  assign n12638_o = n12637_o & n12633_o;
  /* TG68K_ALU.vhd:1202:37  */
  assign n12639_o = result_mulu[63:32];
  /* TG68K_ALU.vhd:1202:51  */
  assign n12641_o = n12639_o == 32'b11111111111111111111111111111111;
  /* TG68K_ALU.vhd:1202:64  */
  assign n12642_o = signedop & n12641_o;
  /* TG68K_ALU.vhd:1202:96  */
  assign n12643_o = result_mulu[31];
  /* TG68K_ALU.vhd:1202:81  */
  assign n12644_o = n12643_o & n12642_o;
  /* TG68K_ALU.vhd:1201:102  */
  assign n12645_o = n12638_o | n12644_o;
  /* TG68K_ALU.vhd:1201:17  */
  assign n12648_o = n12645_o ? 1'b0 : 1'b1;
  /* TG68K_ALU.vhd:1227:77  */
  assign n12653_o = result_mulu[63:32];
  /* TG68K_ALU.vhd:1240:32  */
  assign n12661_o = opcode[15];
  /* TG68K_ALU.vhd:1240:47  */
  assign n12662_o = opcode[8];
  /* TG68K_ALU.vhd:1240:37  */
  assign n12663_o = n12661_o & n12662_o;
  /* TG68K_ALU.vhd:1240:66  */
  assign n12664_o = opcode[15];
  /* TG68K_ALU.vhd:1240:56  */
  assign n12665_o = ~n12664_o;
  /* TG68K_ALU.vhd:1240:81  */
  assign n12666_o = sndopc[11];
  /* TG68K_ALU.vhd:1240:71  */
  assign n12667_o = n12665_o & n12666_o;
  /* TG68K_ALU.vhd:1240:52  */
  assign n12668_o = n12663_o | n12667_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12670_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12671_o = divs & n12670_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12672_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12673_o = divs & n12672_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12674_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12675_o = divs & n12674_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12676_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12677_o = divs & n12676_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12678_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12679_o = divs & n12678_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12680_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12681_o = divs & n12680_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12682_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12683_o = divs & n12682_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12684_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12685_o = divs & n12684_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12686_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12687_o = divs & n12686_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12688_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12689_o = divs & n12688_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12690_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12691_o = divs & n12690_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12692_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12693_o = divs & n12692_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12694_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12695_o = divs & n12694_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12696_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12697_o = divs & n12696_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12698_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12699_o = divs & n12698_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12700_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12701_o = divs & n12700_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12702_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12703_o = divs & n12702_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12704_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12705_o = divs & n12704_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12706_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12707_o = divs & n12706_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12708_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12709_o = divs & n12708_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12710_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12711_o = divs & n12710_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12712_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12713_o = divs & n12712_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12714_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12715_o = divs & n12714_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12716_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12717_o = divs & n12716_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12718_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12719_o = divs & n12718_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12720_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12721_o = divs & n12720_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12722_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12723_o = divs & n12722_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12724_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12725_o = divs & n12724_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12726_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12727_o = divs & n12726_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12728_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12729_o = divs & n12728_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12730_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12731_o = divs & n12730_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12732_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12733_o = divs & n12732_o;
  assign n12734_o = {n12671_o, n12673_o, n12675_o, n12677_o};
  assign n12735_o = {n12679_o, n12681_o, n12683_o, n12685_o};
  assign n12736_o = {n12687_o, n12689_o, n12691_o, n12693_o};
  assign n12737_o = {n12695_o, n12697_o, n12699_o, n12701_o};
  assign n12738_o = {n12703_o, n12705_o, n12707_o, n12709_o};
  assign n12739_o = {n12711_o, n12713_o, n12715_o, n12717_o};
  assign n12740_o = {n12719_o, n12721_o, n12723_o, n12725_o};
  assign n12741_o = {n12727_o, n12729_o, n12731_o, n12733_o};
  assign n12742_o = {n12734_o, n12735_o, n12736_o, n12737_o};
  assign n12743_o = {n12738_o, n12739_o, n12740_o, n12741_o};
  assign n12744_o = {n12742_o, n12743_o};
  /* TG68K_ALU.vhd:1243:30  */
  assign n12745_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1243:39  */
  assign n12747_o = n12745_o | 1'b0;
  /* TG68K_ALU.vhd:1245:52  */
  assign n12748_o = result_div_pre[15];
  /* TG68K_ALU.vhd:1248:38  */
  assign n12749_o = exe_opcode[14];
  /* TG68K_ALU.vhd:1248:57  */
  assign n12750_o = sndopc[10];
  /* TG68K_ALU.vhd:1248:47  */
  assign n12751_o = n12750_o & n12749_o;
  /* TG68K_ALU.vhd:1248:25  */
  assign n12752_o = n12751_o ? reg_qb : n12744_o;
  /* TG68K_ALU.vhd:1251:52  */
  assign n12753_o = result_div_pre[31];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12754_o = n12747_o ? n12748_o : n12753_o;
  assign n12755_o = {n12752_o, reg_qa};
  assign n12756_o = n12755_o[15:0];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12757_o = n12747_o ? 16'b0000000000000000 : n12756_o;
  assign n12758_o = n12755_o[47:16];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12759_o = n12747_o ? reg_qa : n12758_o;
  assign n12760_o = n12755_o[63:48];
  assign n12761_o = n12744_o[31:16];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12762_o = n12747_o ? n12761_o : n12760_o;
  /* TG68K_ALU.vhd:1253:42  */
  assign n12764_o = opcode[15];
  /* TG68K_ALU.vhd:1253:46  */
  assign n12765_o = ~n12764_o;
  /* TG68K_ALU.vhd:1253:33  */
  assign n12766_o = signedop | n12765_o;
  /* TG68K_ALU.vhd:1254:44  */
  assign n12767_o = op2out[31:16];
  /* TG68K_ALU.vhd:1253:17  */
  assign n12769_o = n12766_o ? n12767_o : 16'b0000000000000000;
  /* TG68K_ALU.vhd:1258:43  */
  assign n12770_o = op2out[31];
  /* TG68K_ALU.vhd:1258:33  */
  assign n12771_o = n12770_o & signedop;
  /* TG68K_ALU.vhd:1259:44  */
  assign n12772_o = div_reg[63:31];
  /* TG68K_ALU.vhd:1259:64  */
  assign n12774_o = {1'b1, op2out};
  /* TG68K_ALU.vhd:1259:59  */
  assign n12775_o = n12772_o + n12774_o;
  /* TG68K_ALU.vhd:1261:44  */
  assign n12776_o = div_reg[63:31];
  /* TG68K_ALU.vhd:1261:64  */
  assign n12778_o = {1'b0, op2outext};
  /* TG68K_ALU.vhd:1261:94  */
  assign n12779_o = op2out[15:0];
  /* TG68K_ALU.vhd:1261:87  */
  assign n12780_o = {n12778_o, n12779_o};
  /* TG68K_ALU.vhd:1261:59  */
  assign n12781_o = n12776_o - n12780_o;
  /* TG68K_ALU.vhd:1258:17  */
  assign n12782_o = n12771_o ? n12775_o : n12781_o;
  /* TG68K_ALU.vhd:1266:43  */
  assign n12783_o = div_sub[32];
  /* TG68K_ALU.vhd:1269:58  */
  assign n12784_o = div_reg[62:31];
  /* TG68K_ALU.vhd:1271:58  */
  assign n12785_o = div_sub[31:0];
  /* TG68K_ALU.vhd:1268:17  */
  assign n12786_o = div_bit ? n12784_o : n12785_o;
  /* TG68K_ALU.vhd:1273:49  */
  assign n12787_o = div_reg[30:0];
  /* TG68K_ALU.vhd:1273:63  */
  assign n12788_o = ~div_bit;
  /* TG68K_ALU.vhd:1273:62  */
  assign n12789_o = {n12787_o, n12788_o};
  /* TG68K_ALU.vhd:1276:66  */
  assign n12790_o = div_quot[31:0];
  /* TG68K_ALU.vhd:1276:57  */
  assign n12792_o = 32'b00000000000000000000000000000000 - n12790_o;
  /* TG68K_ALU.vhd:1279:64  */
  assign n12793_o = div_quot[31:0];
  /* TG68K_ALU.vhd:1275:17  */
  assign n12794_o = div_neg ? n12792_o : n12793_o;
  /* TG68K_ALU.vhd:1282:44  */
  assign n12795_o = ~div_bit;
  /* TG68K_ALU.vhd:1282:34  */
  assign n12796_o = nozero | n12795_o;
  /* TG68K_ALU.vhd:1282:50  */
  assign n12797_o = signedop & n12796_o;
  /* TG68K_ALU.vhd:1282:78  */
  assign n12798_o = op2out[31];
  /* TG68K_ALU.vhd:1282:83  */
  assign n12799_o = n12798_o ^ op1_sign;
  /* TG68K_ALU.vhd:1282:96  */
  assign n12800_o = n12799_o ^ div_qsign;
  /* TG68K_ALU.vhd:1282:67  */
  assign n12801_o = n12800_o & n12797_o;
  /* TG68K_ALU.vhd:1283:37  */
  assign n12802_o = ~signedop;
  /* TG68K_ALU.vhd:1283:54  */
  assign n12803_o = div_over[32];
  /* TG68K_ALU.vhd:1283:58  */
  assign n12804_o = ~n12803_o;
  /* TG68K_ALU.vhd:1283:42  */
  assign n12805_o = n12804_o & n12802_o;
  /* TG68K_ALU.vhd:1283:25  */
  assign n12806_o = n12801_o | n12805_o;
  /* TG68K_ALU.vhd:1283:65  */
  assign n12808_o = 1'b1 & n12806_o;
  /* TG68K_ALU.vhd:1282:17  */
  assign n12811_o = n12808_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1294:47  */
  assign n12817_o = micro_state != 7'b1011010;
  /* TG68K_ALU.vhd:1298:47  */
  assign n12820_o = micro_state == 7'b1010101;
  /* TG68K_ALU.vhd:1300:65  */
  assign n12821_o = dividend[63];
  /* TG68K_ALU.vhd:1300:53  */
  assign n12822_o = n12821_o & divs;
  /* TG68K_ALU.vhd:1302:61  */
  assign n12824_o = 64'b0000000000000000000000000000000000000000000000000000000000000000 - dividend;
  /* TG68K_ALU.vhd:1300:41  */
  assign n12825_o = n12822_o ? n12824_o : dividend;
  /* TG68K_ALU.vhd:1300:41  */
  assign n12828_o = n12822_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1309:51  */
  assign n12829_o = ~div_bit;
  /* TG68K_ALU.vhd:1309:63  */
  assign n12830_o = n12829_o | nozero;
  /* TG68K_ALU.vhd:1298:33  */
  assign n12831_o = n12820_o ? n12825_o : div_quot;
  /* TG68K_ALU.vhd:1298:33  */
  assign n12833_o = n12820_o ? 1'b0 : n12830_o;
  /* TG68K_ALU.vhd:1311:47  */
  assign n12836_o = micro_state == 7'b1010110;
  /* TG68K_ALU.vhd:1312:72  */
  assign n12837_o = op2out[31];
  /* TG68K_ALU.vhd:1312:77  */
  assign n12838_o = n12837_o ^ op1_sign;
  /* TG68K_ALU.vhd:1312:61  */
  assign n12839_o = signedop & n12838_o;
  /* TG68K_ALU.vhd:1316:73  */
  assign n12840_o = div_reg[63:32];
  /* TG68K_ALU.vhd:1316:65  */
  assign n12842_o = {1'b0, n12840_o};
  /* TG68K_ALU.vhd:1316:93  */
  assign n12844_o = {1'b0, op2outext};
  /* TG68K_ALU.vhd:1316:123  */
  assign n12845_o = op2out[15:0];
  /* TG68K_ALU.vhd:1316:116  */
  assign n12846_o = {n12844_o, n12845_o};
  /* TG68K_ALU.vhd:1316:88  */
  assign n12847_o = n12842_o - n12846_o;
  /* TG68K_ALU.vhd:1319:40  */
  assign n12850_o = exec[68];
  /* TG68K_ALU.vhd:1319:56  */
  assign n12851_o = ~n12850_o;
  /* TG68K_ALU.vhd:1322:87  */
  assign n12852_o = div_quot[63:32];
  /* TG68K_ALU.vhd:1322:78  */
  assign n12854_o = 32'b00000000000000000000000000000000 - n12852_o;
  /* TG68K_ALU.vhd:1324:85  */
  assign n12855_o = div_quot[63:32];
  /* TG68K_ALU.vhd:1321:41  */
  assign n12856_o = op1_sign ? n12854_o : n12855_o;
  assign n12857_o = {n12856_o, result_div_pre};
  /* TG68K_ALU.vhd:1293:25  */
  assign n12859_o = n12851_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12860_o = n12817_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12862_o = n12836_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12863_o = n12836_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12866_o = n12820_o & clkena_lw;
  assign n12876_o = {n10036_o, n10033_o};
  assign n12877_o = {n10187_o, n10180_o, n10173_o};
  assign n12878_o = {n10165_o, n10164_o, n10159_o, n10117_o};
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12879_q <= n12578_o;
  /* TG68K_ALU.vhd:996:17  */
  assign n12880_o = {n10209_o, n10247_o};
  /* TG68K_ALU.vhd:1292:17  */
  assign n12881_o = n12859_o ? n12857_o : result_div;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12882_q <= n12881_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12883_o = n12860_o ? n12811_o : v_flag;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12884_q <= n12883_o;
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12885_q <= n12579_o;
  /* TG68K_ALU.vhd:405:17  */
  assign n12887_o = clkena_lw ? n10268_o : bchg;
  /* TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n12888_q <= n12887_o;
  /* TG68K_ALU.vhd:405:17  */
  assign n12889_o = clkena_lw ? n10272_o : bset;
  /* TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n12890_q <= n12889_o;
  assign n12894_o = mulu_reg[31:0];
  /* TG68K_ALU.vhd:1211:17  */
  assign n12895_o = clkena_lw ? n12653_o : n12894_o;
  /* TG68K_ALU.vhd:1211:17  */
  always @(posedge clk)
    n12896_q <= n12895_o;
  assign n12898_o = {32'bZ, n12896_q};
  /* TG68K_ALU.vhd:1292:17  */
  assign n12900_o = clkena_lw ? n12831_o : div_reg;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12901_q <= n12900_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12902_o = {n12786_o, n12789_o};
  /* TG68K_ALU.vhd:1292:17  */
  assign n12904_o = n12862_o ? n12839_o : div_neg;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12905_q <= n12904_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12906_o = n12863_o ? n12847_o : div_over;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12907_q <= n12906_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12908_o = clkena_lw ? n12833_o : nozero;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12909_q <= n12908_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12910_o = {n12762_o, n12759_o, n12757_o};
  /* TG68K_ALU.vhd:1292:17  */
  assign n12911_o = clkena_lw ? divs : signedop;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12912_q <= n12911_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12913_o = n12866_o ? n12828_o : op1_sign;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12914_q <= n12913_o;
  assign n12917_o = {n10847_o, n10835_o, n10820_o, n10805_o, n10790_o, n10775_o, n10760_o, n10745_o, n10730_o, n10715_o, n10700_o, n10685_o, n10670_o, n10655_o, n10640_o, n10625_o, n10610_o, n10595_o, n10580_o, n10565_o, n10550_o, n10535_o, n10520_o, n10505_o, n10490_o, n10475_o, n10460_o, n10445_o, n10430_o, n10415_o, n10400_o, n10384_o};
  assign n12919_o = {n11610_o, n11600_o, n11583_o, n11566_o, n11549_o, n11532_o, n11515_o, n11498_o, n11481_o, n11464_o, n11447_o, n11430_o, n11413_o, n11396_o, n11379_o, n11362_o, n11345_o, n11328_o, n11311_o, n11294_o, n11277_o, n11260_o, n11243_o, n11226_o, n11209_o, n11192_o, n11175_o, n11158_o, n11141_o, n11124_o, n11107_o, n11090_o, n11073_o, n11056_o, n11039_o, n11022_o, n11005_o, n10988_o, n10971_o, n10954_o};
  assign n12920_o = {n10848_o, n10840_o, n10825_o, n10810_o, n10795_o, n10780_o, n10765_o, n10750_o, n10735_o, n10720_o, n10705_o, n10690_o, n10675_o, n10660_o, n10645_o, n10630_o, n10615_o, n10600_o, n10585_o, n10570_o, n10555_o, n10540_o, n10525_o, n10510_o, n10495_o, n10480_o, n10465_o, n10450_o, n10435_o, n10420_o, n10405_o, n10389_o};
  assign n12922_o = {n10904_o, n10905_o};
  assign n12923_o = {n11694_o, n11723_o, n11720_o};
  /* TG68K_ALU.vhd:446:17  */
  assign n12924_o = clkena_lw ? n10331_o : bf_bset;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12925_q <= n12924_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12926_o = clkena_lw ? n10335_o : bf_bchg;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12927_q <= n12926_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12928_o = clkena_lw ? n10339_o : bf_ins;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12929_q <= n12928_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12930_o = clkena_lw ? n10343_o : bf_exts;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12931_q <= n12930_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12932_o = clkena_lw ? n10347_o : bf_fffo;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12933_q <= n12932_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12934_o = clkena_lw ? n10356_o : bf_d32;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12935_q <= n12934_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12936_o = clkena_lw ? n10350_o : bf_s32;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12937_q <= n12936_o;
  assign n12939_o = {n12214_o, n12212_o, n12209_o, n12206_o, n12203_o, n12216_o};
  assign n12940_o = {n11895_o, n11892_o, n11896_o, n11890_o, n11894_o};
  assign n12941_o = {n12149_o, n12151_o};
  assign n12942_o = {n12230_o, n12225_o, n12236_o};
  /* TG68K_ALU.vhd:446:17  */
  assign n12943_o = clkena_lw ? n10358_o : n12944_q;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12944_q <= n12943_o;
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12945_q <= n12586_o;
  /* TG68K_ALU.vhd:76:17  */
  assign n12946_o = op1out[0];
  /* TG68K_ALU.vhd:75:17  */
  assign n12947_o = op1out[1];
  /* TG68K_ALU.vhd:74:17  */
  assign n12948_o = op1out[2];
  /* TG68K_ALU.vhd:73:17  */
  assign n12949_o = op1out[3];
  /* TG68K_ALU.vhd:72:17  */
  assign n12950_o = op1out[4];
  /* TG68K_ALU.vhd:66:17  */
  assign n12951_o = op1out[5];
  /* TG68K_ALU.vhd:446:17  */
  assign n12952_o = op1out[6];
  assign n12953_o = op1out[7];
  assign n12954_o = op1out[8];
  assign n12955_o = op1out[9];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12956_o = op1out[10];
  assign n12957_o = op1out[11];
  assign n12958_o = op1out[12];
  assign n12959_o = op1out[13];
  assign n12960_o = op1out[14];
  /* TG68K_ALU.vhd:405:17  */
  assign n12961_o = op1out[15];
  /* TG68K_ALU.vhd:996:17  */
  assign n12962_o = op1out[16];
  assign n12963_o = op1out[17];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12964_o = op1out[18];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12965_o = op1out[19];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12966_o = op1out[20];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12967_o = op1out[21];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12968_o = op1out[22];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12969_o = op1out[23];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12970_o = op1out[24];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12971_o = op1out[25];
  /* TG68K_ALU.vhd:1290:1  */
  assign n12972_o = op1out[26];
  assign n12973_o = op1out[27];
  assign n12974_o = op1out[28];
  /* TG68K_ALU.vhd:1237:1  */
  assign n12975_o = op1out[29];
  assign n12976_o = op1out[30];
  /* TG68K_ALU.vhd:1211:17  */
  assign n12977_o = op1out[31];
  /* TG68K_ALU.vhd:433:37  */
  assign n12978_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12978_o)
      2'b00: n12979_o = n12946_o;
      2'b01: n12979_o = n12947_o;
      2'b10: n12979_o = n12948_o;
      2'b11: n12979_o = n12949_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12980_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12980_o)
      2'b00: n12981_o = n12950_o;
      2'b01: n12981_o = n12951_o;
      2'b10: n12981_o = n12952_o;
      2'b11: n12981_o = n12953_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12982_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12982_o)
      2'b00: n12983_o = n12954_o;
      2'b01: n12983_o = n12955_o;
      2'b10: n12983_o = n12956_o;
      2'b11: n12983_o = n12957_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12984_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12984_o)
      2'b00: n12985_o = n12958_o;
      2'b01: n12985_o = n12959_o;
      2'b10: n12985_o = n12960_o;
      2'b11: n12985_o = n12961_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12986_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12986_o)
      2'b00: n12987_o = n12962_o;
      2'b01: n12987_o = n12963_o;
      2'b10: n12987_o = n12964_o;
      2'b11: n12987_o = n12965_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12988_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12988_o)
      2'b00: n12989_o = n12966_o;
      2'b01: n12989_o = n12967_o;
      2'b10: n12989_o = n12968_o;
      2'b11: n12989_o = n12969_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12990_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12990_o)
      2'b00: n12991_o = n12970_o;
      2'b01: n12991_o = n12971_o;
      2'b10: n12991_o = n12972_o;
      2'b11: n12991_o = n12973_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12992_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12992_o)
      2'b00: n12993_o = n12974_o;
      2'b01: n12993_o = n12975_o;
      2'b10: n12993_o = n12976_o;
      2'b11: n12993_o = n12977_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12994_o = bit_number[3:2];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12994_o)
      2'b00: n12995_o = n12979_o;
      2'b01: n12995_o = n12981_o;
      2'b10: n12995_o = n12983_o;
      2'b11: n12995_o = n12985_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12996_o = bit_number[3:2];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12996_o)
      2'b00: n12997_o = n12987_o;
      2'b01: n12997_o = n12989_o;
      2'b10: n12997_o = n12991_o;
      2'b11: n12997_o = n12993_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12998_o = bit_number[4];
  /* TG68K_ALU.vhd:433:37  */
  assign n12999_o = n12998_o ? n12997_o : n12995_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13000_o = bit_number[4];
  /* TG68K_ALU.vhd:435:17  */
  assign n13001_o = ~n13000_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13002_o = bit_number[3];
  /* TG68K_ALU.vhd:435:17  */
  assign n13003_o = ~n13002_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13004_o = n13001_o & n13003_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13005_o = n13001_o & n13002_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13006_o = n13000_o & n13003_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13007_o = n13000_o & n13002_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13008_o = bit_number[2];
  /* TG68K_ALU.vhd:435:17  */
  assign n13009_o = ~n13008_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13010_o = n13004_o & n13009_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13011_o = n13004_o & n13008_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13012_o = n13005_o & n13009_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13013_o = n13005_o & n13008_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13014_o = n13006_o & n13009_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13015_o = n13006_o & n13008_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13016_o = n13007_o & n13009_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13017_o = n13007_o & n13008_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13018_o = bit_number[1];
  /* TG68K_ALU.vhd:435:17  */
  assign n13019_o = ~n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13020_o = n13010_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13021_o = n13010_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13022_o = n13011_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13023_o = n13011_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13024_o = n13012_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13025_o = n13012_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13026_o = n13013_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13027_o = n13013_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13028_o = n13014_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13029_o = n13014_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13030_o = n13015_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13031_o = n13015_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13032_o = n13016_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13033_o = n13016_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13034_o = n13017_o & n13019_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13035_o = n13017_o & n13018_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13036_o = bit_number[0];
  /* TG68K_ALU.vhd:435:17  */
  assign n13037_o = ~n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13038_o = n13020_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13039_o = n13020_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13040_o = n13021_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13041_o = n13021_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13042_o = n13022_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13043_o = n13022_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13044_o = n13023_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13045_o = n13023_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13046_o = n13024_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13047_o = n13024_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13048_o = n13025_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13049_o = n13025_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13050_o = n13026_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13051_o = n13026_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13052_o = n13027_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13053_o = n13027_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13054_o = n13028_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13055_o = n13028_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13056_o = n13029_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13057_o = n13029_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13058_o = n13030_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13059_o = n13030_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13060_o = n13031_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13061_o = n13031_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13062_o = n13032_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13063_o = n13032_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13064_o = n13033_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13065_o = n13033_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13066_o = n13034_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13067_o = n13034_o & n13036_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13068_o = n13035_o & n13037_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n13069_o = n13035_o & n13036_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13070_o = op1out[0];
  /* TG68K_ALU.vhd:435:17  */
  assign n13071_o = n13038_o ? n10304_o : n13070_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13072_o = op1out[1];
  /* TG68K_ALU.vhd:435:17  */
  assign n13073_o = n13039_o ? n10304_o : n13072_o;
  assign n13074_o = op1out[2];
  /* TG68K_ALU.vhd:435:17  */
  assign n13075_o = n13040_o ? n10304_o : n13074_o;
  assign n13076_o = op1out[3];
  /* TG68K_ALU.vhd:435:17  */
  assign n13077_o = n13041_o ? n10304_o : n13076_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13078_o = op1out[4];
  /* TG68K_ALU.vhd:435:17  */
  assign n13079_o = n13042_o ? n10304_o : n13078_o;
  assign n13080_o = op1out[5];
  /* TG68K_ALU.vhd:435:17  */
  assign n13081_o = n13043_o ? n10304_o : n13080_o;
  assign n13082_o = op1out[6];
  /* TG68K_ALU.vhd:435:17  */
  assign n13083_o = n13044_o ? n10304_o : n13082_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13084_o = op1out[7];
  /* TG68K_ALU.vhd:435:17  */
  assign n13085_o = n13045_o ? n10304_o : n13084_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13086_o = op1out[8];
  /* TG68K_ALU.vhd:435:17  */
  assign n13087_o = n13046_o ? n10304_o : n13086_o;
  assign n13088_o = op1out[9];
  /* TG68K_ALU.vhd:435:17  */
  assign n13089_o = n13047_o ? n10304_o : n13088_o;
  assign n13090_o = op1out[10];
  /* TG68K_ALU.vhd:435:17  */
  assign n13091_o = n13048_o ? n10304_o : n13090_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13092_o = op1out[11];
  /* TG68K_ALU.vhd:435:17  */
  assign n13093_o = n13049_o ? n10304_o : n13092_o;
  assign n13094_o = op1out[12];
  /* TG68K_ALU.vhd:435:17  */
  assign n13095_o = n13050_o ? n10304_o : n13094_o;
  assign n13096_o = op1out[13];
  /* TG68K_ALU.vhd:435:17  */
  assign n13097_o = n13051_o ? n10304_o : n13096_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13098_o = op1out[14];
  /* TG68K_ALU.vhd:435:17  */
  assign n13099_o = n13052_o ? n10304_o : n13098_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13100_o = op1out[15];
  /* TG68K_ALU.vhd:435:17  */
  assign n13101_o = n13053_o ? n10304_o : n13100_o;
  assign n13102_o = op1out[16];
  /* TG68K_ALU.vhd:435:17  */
  assign n13103_o = n13054_o ? n10304_o : n13102_o;
  assign n13104_o = op1out[17];
  /* TG68K_ALU.vhd:435:17  */
  assign n13105_o = n13055_o ? n10304_o : n13104_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13106_o = op1out[18];
  /* TG68K_ALU.vhd:435:17  */
  assign n13107_o = n13056_o ? n10304_o : n13106_o;
  assign n13108_o = op1out[19];
  /* TG68K_ALU.vhd:435:17  */
  assign n13109_o = n13057_o ? n10304_o : n13108_o;
  assign n13110_o = op1out[20];
  /* TG68K_ALU.vhd:435:17  */
  assign n13111_o = n13058_o ? n10304_o : n13110_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13112_o = op1out[21];
  /* TG68K_ALU.vhd:435:17  */
  assign n13113_o = n13059_o ? n10304_o : n13112_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13114_o = op1out[22];
  /* TG68K_ALU.vhd:435:17  */
  assign n13115_o = n13060_o ? n10304_o : n13114_o;
  assign n13116_o = op1out[23];
  /* TG68K_ALU.vhd:435:17  */
  assign n13117_o = n13061_o ? n10304_o : n13116_o;
  assign n13118_o = op1out[24];
  /* TG68K_ALU.vhd:435:17  */
  assign n13119_o = n13062_o ? n10304_o : n13118_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13120_o = op1out[25];
  /* TG68K_ALU.vhd:435:17  */
  assign n13121_o = n13063_o ? n10304_o : n13120_o;
  assign n13122_o = op1out[26];
  /* TG68K_ALU.vhd:435:17  */
  assign n13123_o = n13064_o ? n10304_o : n13122_o;
  assign n13124_o = op1out[27];
  /* TG68K_ALU.vhd:435:17  */
  assign n13125_o = n13065_o ? n10304_o : n13124_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13126_o = op1out[28];
  /* TG68K_ALU.vhd:435:17  */
  assign n13127_o = n13066_o ? n10304_o : n13126_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13128_o = op1out[29];
  /* TG68K_ALU.vhd:435:17  */
  assign n13129_o = n13067_o ? n10304_o : n13128_o;
  assign n13130_o = op1out[30];
  /* TG68K_ALU.vhd:435:17  */
  assign n13131_o = n13068_o ? n10304_o : n13130_o;
  assign n13132_o = op1out[31];
  /* TG68K_ALU.vhd:435:17  */
  assign n13133_o = n13069_o ? n10304_o : n13132_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13134_o = {n13133_o, n13131_o, n13129_o, n13127_o, n13125_o, n13123_o, n13121_o, n13119_o, n13117_o, n13115_o, n13113_o, n13111_o, n13109_o, n13107_o, n13105_o, n13103_o, n13101_o, n13099_o, n13097_o, n13095_o, n13093_o, n13091_o, n13089_o, n13087_o, n13085_o, n13083_o, n13081_o, n13079_o, n13077_o, n13075_o, n13073_o, n13071_o};
  /* TG68K_ALU.vhd:435:26  */
  assign n13135_o = datareg[0];
  /* TG68K_ALU.vhd:435:17  */
  assign n13136_o = datareg[1];
  /* TG68K_ALU.vhd:575:17  */
  assign n13137_o = datareg[2];
  assign n13138_o = datareg[3];
  assign n13139_o = datareg[4];
  assign n13140_o = datareg[5];
  assign n13141_o = datareg[6];
  /* TG68K_ALU.vhd:581:17  */
  assign n13142_o = datareg[7];
  /* TG68K_ALU.vhd:572:17  */
  assign n13143_o = datareg[8];
  /* TG68K_ALU.vhd:575:17  */
  assign n13144_o = datareg[9];
  assign n13145_o = datareg[10];
  assign n13146_o = datareg[11];
  assign n13147_o = datareg[12];
  assign n13148_o = datareg[13];
  /* TG68K_ALU.vhd:581:17  */
  assign n13149_o = datareg[14];
  /* TG68K_ALU.vhd:572:17  */
  assign n13150_o = datareg[15];
  /* TG68K_ALU.vhd:575:17  */
  assign n13151_o = datareg[16];
  assign n13152_o = datareg[17];
  assign n13153_o = datareg[18];
  assign n13154_o = datareg[19];
  assign n13155_o = datareg[20];
  /* TG68K_ALU.vhd:581:17  */
  assign n13156_o = datareg[21];
  /* TG68K_ALU.vhd:572:17  */
  assign n13157_o = datareg[22];
  /* TG68K_ALU.vhd:575:17  */
  assign n13158_o = datareg[23];
  assign n13159_o = datareg[24];
  assign n13160_o = datareg[25];
  assign n13161_o = datareg[26];
  assign n13162_o = datareg[27];
  /* TG68K_ALU.vhd:581:17  */
  assign n13163_o = datareg[28];
  /* TG68K_ALU.vhd:572:17  */
  assign n13164_o = datareg[29];
  /* TG68K_ALU.vhd:575:17  */
  assign n13165_o = datareg[30];
  assign n13166_o = datareg[31];
  /* TG68K_ALU.vhd:496:36  */
  assign n13167_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13167_o)
      2'b00: n13168_o = n13135_o;
      2'b01: n13168_o = n13136_o;
      2'b10: n13168_o = n13137_o;
      2'b11: n13168_o = n13138_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13169_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13169_o)
      2'b00: n13170_o = n13139_o;
      2'b01: n13170_o = n13140_o;
      2'b10: n13170_o = n13141_o;
      2'b11: n13170_o = n13142_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13171_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13171_o)
      2'b00: n13172_o = n13143_o;
      2'b01: n13172_o = n13144_o;
      2'b10: n13172_o = n13145_o;
      2'b11: n13172_o = n13146_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13173_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13173_o)
      2'b00: n13174_o = n13147_o;
      2'b01: n13174_o = n13148_o;
      2'b10: n13174_o = n13149_o;
      2'b11: n13174_o = n13150_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13175_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13175_o)
      2'b00: n13176_o = n13151_o;
      2'b01: n13176_o = n13152_o;
      2'b10: n13176_o = n13153_o;
      2'b11: n13176_o = n13154_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13177_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13177_o)
      2'b00: n13178_o = n13155_o;
      2'b01: n13178_o = n13156_o;
      2'b10: n13178_o = n13157_o;
      2'b11: n13178_o = n13158_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13179_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13179_o)
      2'b00: n13180_o = n13159_o;
      2'b01: n13180_o = n13160_o;
      2'b10: n13180_o = n13161_o;
      2'b11: n13180_o = n13162_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13181_o = n10850_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13181_o)
      2'b00: n13182_o = n13163_o;
      2'b01: n13182_o = n13164_o;
      2'b10: n13182_o = n13165_o;
      2'b11: n13182_o = n13166_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13183_o = n10850_o[3:2];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13183_o)
      2'b00: n13184_o = n13168_o;
      2'b01: n13184_o = n13170_o;
      2'b10: n13184_o = n13172_o;
      2'b11: n13184_o = n13174_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13185_o = n10850_o[3:2];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13185_o)
      2'b00: n13186_o = n13176_o;
      2'b01: n13186_o = n13178_o;
      2'b10: n13186_o = n13180_o;
      2'b11: n13186_o = n13182_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13187_o = n10850_o[4];
  /* TG68K_ALU.vhd:496:36  */
  assign n13188_o = n13187_o ? n13186_o : n13184_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13189_o = bit_msb[5];
  /* TG68K_ALU.vhd:761:17  */
  assign n13190_o = ~n13189_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13191_o = bit_msb[4];
  /* TG68K_ALU.vhd:761:17  */
  assign n13192_o = ~n13191_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13193_o = n13190_o & n13192_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13194_o = n13190_o & n13191_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13195_o = n13189_o & n13192_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13196_o = bit_msb[3];
  /* TG68K_ALU.vhd:761:17  */
  assign n13197_o = ~n13196_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13198_o = n13193_o & n13197_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13199_o = n13193_o & n13196_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13200_o = n13194_o & n13197_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13201_o = n13194_o & n13196_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13202_o = n13195_o & n13197_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13203_o = bit_msb[2];
  /* TG68K_ALU.vhd:761:17  */
  assign n13204_o = ~n13203_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13205_o = n13198_o & n13204_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13206_o = n13198_o & n13203_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13207_o = n13199_o & n13204_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13208_o = n13199_o & n13203_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13209_o = n13200_o & n13204_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13210_o = n13200_o & n13203_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13211_o = n13201_o & n13204_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13212_o = n13201_o & n13203_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13213_o = n13202_o & n13204_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13214_o = bit_msb[1];
  /* TG68K_ALU.vhd:761:17  */
  assign n13215_o = ~n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13216_o = n13205_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13217_o = n13205_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13218_o = n13206_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13219_o = n13206_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13220_o = n13207_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13221_o = n13207_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13222_o = n13208_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13223_o = n13208_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13224_o = n13209_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13225_o = n13209_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13226_o = n13210_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13227_o = n13210_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13228_o = n13211_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13229_o = n13211_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13230_o = n13212_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13231_o = n13212_o & n13214_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13232_o = n13213_o & n13215_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13233_o = bit_msb[0];
  /* TG68K_ALU.vhd:761:17  */
  assign n13234_o = ~n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13235_o = n13216_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13236_o = n13216_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13237_o = n13217_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13238_o = n13217_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13239_o = n13218_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13240_o = n13218_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13241_o = n13219_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13242_o = n13219_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13243_o = n13220_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13244_o = n13220_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13245_o = n13221_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13246_o = n13221_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13247_o = n13222_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13248_o = n13222_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13249_o = n13223_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13250_o = n13223_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13251_o = n13224_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13252_o = n13224_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13253_o = n13225_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13254_o = n13225_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13255_o = n13226_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13256_o = n13226_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13257_o = n13227_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13258_o = n13227_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13259_o = n13228_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13260_o = n13228_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13261_o = n13229_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13262_o = n13229_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13263_o = n13230_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13264_o = n13230_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13265_o = n13231_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13266_o = n13231_o & n13233_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13267_o = n13232_o & n13234_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13268_o = n13232_o & n13233_o;
  assign n13269_o = n11861_o[0];
  /* TG68K_ALU.vhd:761:17  */
  assign n13270_o = n13235_o ? 1'b1 : n13269_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13271_o = n11861_o[1];
  /* TG68K_ALU.vhd:761:17  */
  assign n13272_o = n13236_o ? 1'b1 : n13271_o;
  assign n13273_o = n11861_o[2];
  /* TG68K_ALU.vhd:761:17  */
  assign n13274_o = n13237_o ? 1'b1 : n13273_o;
  assign n13275_o = n11861_o[3];
  /* TG68K_ALU.vhd:761:17  */
  assign n13276_o = n13238_o ? 1'b1 : n13275_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13277_o = n11861_o[4];
  /* TG68K_ALU.vhd:761:17  */
  assign n13278_o = n13239_o ? 1'b1 : n13277_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13279_o = n11861_o[5];
  /* TG68K_ALU.vhd:761:17  */
  assign n13280_o = n13240_o ? 1'b1 : n13279_o;
  assign n13281_o = n11861_o[6];
  /* TG68K_ALU.vhd:761:17  */
  assign n13282_o = n13241_o ? 1'b1 : n13281_o;
  assign n13283_o = n11861_o[7];
  /* TG68K_ALU.vhd:761:17  */
  assign n13284_o = n13242_o ? 1'b1 : n13283_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13285_o = n11861_o[8];
  /* TG68K_ALU.vhd:761:17  */
  assign n13286_o = n13243_o ? 1'b1 : n13285_o;
  assign n13287_o = n11861_o[9];
  /* TG68K_ALU.vhd:761:17  */
  assign n13288_o = n13244_o ? 1'b1 : n13287_o;
  assign n13289_o = n11861_o[10];
  /* TG68K_ALU.vhd:761:17  */
  assign n13290_o = n13245_o ? 1'b1 : n13289_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13291_o = n11861_o[11];
  /* TG68K_ALU.vhd:761:17  */
  assign n13292_o = n13246_o ? 1'b1 : n13291_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13293_o = n11861_o[12];
  /* TG68K_ALU.vhd:761:17  */
  assign n13294_o = n13247_o ? 1'b1 : n13293_o;
  assign n13295_o = n11861_o[13];
  /* TG68K_ALU.vhd:761:17  */
  assign n13296_o = n13248_o ? 1'b1 : n13295_o;
  assign n13297_o = n11861_o[14];
  /* TG68K_ALU.vhd:761:17  */
  assign n13298_o = n13249_o ? 1'b1 : n13297_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13299_o = n11861_o[15];
  /* TG68K_ALU.vhd:761:17  */
  assign n13300_o = n13250_o ? 1'b1 : n13299_o;
  assign n13301_o = n11861_o[16];
  /* TG68K_ALU.vhd:761:17  */
  assign n13302_o = n13251_o ? 1'b1 : n13301_o;
  assign n13303_o = n11861_o[17];
  /* TG68K_ALU.vhd:761:17  */
  assign n13304_o = n13252_o ? 1'b1 : n13303_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13305_o = n11861_o[18];
  /* TG68K_ALU.vhd:761:17  */
  assign n13306_o = n13253_o ? 1'b1 : n13305_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13307_o = n11861_o[19];
  /* TG68K_ALU.vhd:761:17  */
  assign n13308_o = n13254_o ? 1'b1 : n13307_o;
  assign n13309_o = n11861_o[20];
  /* TG68K_ALU.vhd:761:17  */
  assign n13310_o = n13255_o ? 1'b1 : n13309_o;
  assign n13311_o = n11861_o[21];
  /* TG68K_ALU.vhd:761:17  */
  assign n13312_o = n13256_o ? 1'b1 : n13311_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13313_o = n11861_o[22];
  /* TG68K_ALU.vhd:761:17  */
  assign n13314_o = n13257_o ? 1'b1 : n13313_o;
  assign n13315_o = n11861_o[23];
  /* TG68K_ALU.vhd:761:17  */
  assign n13316_o = n13258_o ? 1'b1 : n13315_o;
  assign n13317_o = n11861_o[24];
  /* TG68K_ALU.vhd:761:17  */
  assign n13318_o = n13259_o ? 1'b1 : n13317_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13319_o = n11861_o[25];
  /* TG68K_ALU.vhd:761:17  */
  assign n13320_o = n13260_o ? 1'b1 : n13319_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13321_o = n11861_o[26];
  /* TG68K_ALU.vhd:761:17  */
  assign n13322_o = n13261_o ? 1'b1 : n13321_o;
  assign n13323_o = n11861_o[27];
  /* TG68K_ALU.vhd:761:17  */
  assign n13324_o = n13262_o ? 1'b1 : n13323_o;
  assign n13325_o = n11861_o[28];
  /* TG68K_ALU.vhd:761:17  */
  assign n13326_o = n13263_o ? 1'b1 : n13325_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13327_o = n11861_o[29];
  /* TG68K_ALU.vhd:761:17  */
  assign n13328_o = n13264_o ? 1'b1 : n13327_o;
  assign n13329_o = n11861_o[30];
  /* TG68K_ALU.vhd:761:17  */
  assign n13330_o = n13265_o ? 1'b1 : n13329_o;
  assign n13331_o = n11861_o[31];
  /* TG68K_ALU.vhd:761:17  */
  assign n13332_o = n13266_o ? 1'b1 : n13331_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13333_o = n11861_o[32];
  /* TG68K_ALU.vhd:761:17  */
  assign n13334_o = n13267_o ? 1'b1 : n13333_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13335_o = n11861_o[33];
  /* TG68K_ALU.vhd:761:17  */
  assign n13336_o = n13268_o ? 1'b1 : n13335_o;
  assign n13337_o = {n13336_o, n13334_o, n13332_o, n13330_o, n13328_o, n13326_o, n13324_o, n13322_o, n13320_o, n13318_o, n13316_o, n13314_o, n13312_o, n13310_o, n13308_o, n13306_o, n13304_o, n13302_o, n13300_o, n13298_o, n13296_o, n13294_o, n13292_o, n13290_o, n13288_o, n13286_o, n13284_o, n13282_o, n13280_o, n13278_o, n13276_o, n13274_o, n13272_o, n13270_o};
endmodule

module tg68kdotc_kernel_2_2_2_2_2_2_1_1
  (input  clk,
   input  nreset,
   input  clkena_in,
   input  [15:0] data_in,
   input  [2:0] ipl,
   input  ipl_autovector,
   input  berr,
   input  [1:0] cpu,
   output [31:0] addr_out,
   output [15:0] data_write,
   output nwr,
   output nuds,
   output nlds,
   output [1:0] busstate,
   output longword,
   output nresetout,
   output [2:0] fc,
   output clr_berr,
   output skipfetch,
   output [31:0] regin_out,
   output [3:0] cacr_out,
   output [31:0] vbr_out);
  wire use_vbr_stackframe;
  wire [3:0] syncreset;
  wire reset;
  wire clkena_lw;
  wire [31:0] tg68_pc;
  wire [31:0] tmp_tg68_pc;
  wire [31:0] tg68_pc_add;
  wire [31:0] pc_dataa;
  wire [31:0] pc_datab;
  wire [31:0] memaddr;
  wire [1:0] state;
  wire [1:0] datatype;
  wire [1:0] set_datatype;
  wire [1:0] exe_datatype;
  wire [1:0] setstate;
  wire setaddrvalue;
  wire addrvalue;
  wire [15:0] opcode;
  wire [15:0] exe_opcode;
  wire [15:0] sndopc;
  wire [31:0] exe_pc  /*verilator public_flat_rd*/ ;
  wire [31:0] last_opc_pc;
  wire [15:0] last_opc_read;
  wire [31:0] reg_qa;
  wire [31:0] reg_qb;
  wire wwrena;
  wire lwrena;
  wire bwrena;
  wire regwrena_now;
  wire [3:0] rf_dest_addr;
  wire [3:0] rf_source_addr;
  wire [3:0] rf_source_addrd;
  wire [31:0] regin;
  wire [3:0] rdindex_a;
  wire [3:0] rdindex_b;
  wire wr_areg;
  wire [31:0] addr;
  wire [31:0] memaddr_reg;
  wire [31:0] memaddr_delta;
  wire [31:0] memaddr_delta_rega;
  wire [31:0] memaddr_delta_regb;
  wire use_base;
  wire [31:0] ea_data;
  wire [31:0] op1out;
  wire [31:0] op2out;
  wire [15:0] op1outbrief;
  wire [31:0] aluout;
  wire [31:0] data_write_tmp;
  wire [31:0] data_write_muxin;
  wire [47:0] data_write_mux;
  wire nextpass;
  wire setnextpass;
  wire setdispbyte;
  wire setdisp;
  wire regdirectsource;
  wire [31:0] addsub_q;
  wire [31:0] briefdata;
  wire [2:0] c_out;
  wire [31:0] memaddr_a;
  wire tg68_pc_brw;
  wire tg68_pc_word;
  wire getbrief;
  wire [15:0] brief;
  wire data_is_source;
  wire store_in_tmp;
  wire write_back;
  wire exec_write_back;
  wire setstackaddr;
  wire writepc;
  wire writepcbig;
  wire set_writepcbig;
  wire writepcnext;
  wire setopcode;
  wire decodeopc  /*verilator public_flat_rd*/ ;
  wire execopc;
  wire execopc_alu;
  wire setexecopc;
  wire endopc;
  wire setendopc;
  wire [7:0] flags;
  wire [7:0] flagssr;
  wire [7:0] srin;
  wire exec_direct;
  wire exec_tas;
  wire set_exec_tas;
  wire exe_condition;
  wire ea_only;
  wire source_areg;
  wire source_lowbits;
  wire source_ldrlbits;
  wire source_ldrmbits;
  wire source_2ndhbits;
  wire source_2ndmbits;
  wire source_2ndlbits;
  wire dest_areg;
  wire dest_ldrareg;
  wire dest_ldrhbits;
  wire dest_ldrlbits;
  wire dest_2ndhbits;
  wire dest_2ndlbits;
  wire dest_hbits;
  wire [1:0] rot_bits;
  wire [1:0] set_rot_bits;
  wire [5:0] rot_cnt;
  wire [5:0] set_rot_cnt;
  wire movem_actiond;
  wire [3:0] movem_regaddr;
  wire [3:0] movem_mux;
  wire movem_presub;
  wire movem_run;
  wire set_direct_data;
  wire use_direct_data;
  wire direct_data;
  wire set_v_flag;
  wire set_vectoraddr;
  wire writesr;
  wire trap_berr;
  wire trap_illegal;
  wire trap_addr_error;
  wire trap_priv;
  wire trap_trace;
  wire trap_1010;
  wire trap_1111;
  wire trap_trap;
  wire trap_trapv;
  wire trap_interrupt;
  wire trapmake;
  wire trapd;
  wire [7:0] trap_sr;
  wire make_trace;
  wire make_berr;
  wire usestackframe2;
  wire set_stop;
  wire stop;
  wire [31:0] trap_vector;
  wire [31:0] trap_vector_vbr;
  wire [31:0] usp;
  wire [2:0] ipl_nr;
  wire [2:0] ripl_nr;
  wire [7:0] ipl_vec;
  wire interrupt;
  wire setinterrupt;
  wire svmode;
  wire presvmode;
  wire suppress_base;
  wire set_suppress_base;
  wire set_z_error;
  wire z_error;
  wire ea_build_now;
  wire build_logical;
  wire build_bcd;
  wire [31:0] data_read;
  wire [7:0] bf_ext_in;
  wire [7:0] bf_ext_out;
  wire long_start;
  wire long_start_alu;
  wire non_aligned;
  wire check_aligned;
  wire long_done;
  wire [5:0] memmask;
  wire [5:0] set_memmask;
  wire [3:0] memread;
  wire [5:0] wbmemmask;
  wire [5:0] memmaskmux;
  wire oddout;
  wire set_oddout;
  wire pcbase;
  wire set_pcbase;
  wire [31:0] last_data_read;
  wire [31:0] last_data_in;
  wire [5:0] bf_offset;
  wire [5:0] bf_width;
  wire [5:0] bf_bhits;
  wire [5:0] bf_shift;
  wire [5:0] alu_width;
  wire [5:0] alu_bf_shift;
  wire [5:0] bf_loffset;
  wire [31:0] bf_full_offset;
  wire [31:0] alu_bf_ffo_offset;
  wire [5:0] alu_bf_loffset;
  wire [31:0] movec_data;
  wire [31:0] vbr;
  wire [3:0] cacr;
  wire [2:0] dfc;
  wire [2:0] sfc;
  wire [88:0] set;
  wire [88:0] set_exec;
  wire [88:0] exec;
  wire [6:0] micro_state;
  wire [6:0] next_micro_state;
  wire [15:0] n34_o;
  wire [15:0] n35_o;
  wire [7:0] alu_n36;
  wire [4:0] n37_o;
  wire alu_n38;
  wire [7:0] alu_n39;
  wire [2:0] alu_n40;
  wire [31:0] alu_n41;
  wire [31:0] alu_n42;
  wire [7:0] alu_bf_ext_out;
  wire alu_set_v_flag;
  wire [7:0] alu_flags;
  wire [2:0] alu_c_out;
  wire [31:0] alu_addsub_q;
  wire [31:0] alu_aluout;
  wire n55_o;
  wire n56_o;
  wire n57_o;
  wire n58_o;
  wire n59_o;
  wire n60_o;
  wire [1:0] n63_o;
  wire n65_o;
  wire [1:0] n66_o;
  wire n68_o;
  wire n69_o;
  wire n72_o;
  wire n77_o;
  wire n78_o;
  wire n81_o;
  wire n82_o;
  wire n84_o;
  wire [5:0] n85_o;
  wire [4:0] n86_o;
  wire [5:0] n88_o;
  wire n89_o;
  wire n90_o;
  wire n92_o;
  wire n93_o;
  wire n94_o;
  wire n97_o;
  wire n98_o;
  wire n102_o;
  wire [2:0] n104_o;
  wire [3:0] n106_o;
  wire n107_o;
  wire n108_o;
  wire n118_o;
  wire n120_o;
  wire n122_o;
  wire n125_o;
  wire n130_o;
  wire n131_o;
  wire [15:0] n132_o;
  wire [31:0] n133_o;
  wire [23:0] n134_o;
  wire [7:0] n135_o;
  wire [31:0] n136_o;
  wire n138_o;
  wire [1:0] n139_o;
  wire n141_o;
  wire n142_o;
  wire n143_o;
  wire n144_o;
  wire n145_o;
  wire n146_o;
  wire n147_o;
  wire n148_o;
  wire n149_o;
  wire n150_o;
  wire n151_o;
  wire n152_o;
  wire n153_o;
  wire n154_o;
  wire n155_o;
  wire n156_o;
  wire n157_o;
  wire n158_o;
  wire n159_o;
  wire n160_o;
  wire [3:0] n161_o;
  wire [3:0] n162_o;
  wire [3:0] n163_o;
  wire [3:0] n164_o;
  wire [15:0] n165_o;
  wire [15:0] n166_o;
  wire [15:0] n167_o;
  wire [15:0] n168_o;
  wire [15:0] n169_o;
  wire [15:0] n170_o;
  wire [15:0] n171_o;
  wire [15:0] n172_o;
  wire n175_o;
  wire n176_o;
  wire n177_o;
  wire n178_o;
  wire [7:0] n179_o;
  wire [7:0] n180_o;
  wire [7:0] n181_o;
  wire n184_o;
  wire n185_o;
  wire n186_o;
  wire n187_o;
  wire n188_o;
  wire n189_o;
  wire n190_o;
  wire n191_o;
  wire n192_o;
  wire n193_o;
  wire n194_o;
  wire n195_o;
  wire n196_o;
  wire n197_o;
  wire n198_o;
  wire n199_o;
  wire n200_o;
  wire n201_o;
  wire n202_o;
  wire n203_o;
  wire n204_o;
  wire n205_o;
  wire n206_o;
  wire n207_o;
  wire n208_o;
  wire n209_o;
  wire n210_o;
  wire n211_o;
  wire [3:0] n212_o;
  wire [3:0] n213_o;
  wire [3:0] n214_o;
  wire [3:0] n215_o;
  wire [15:0] n216_o;
  wire [15:0] n217_o;
  wire [15:0] n218_o;
  wire [15:0] n219_o;
  wire [15:0] n220_o;
  wire [31:0] n221_o;
  wire [31:0] n222_o;
  wire [15:0] n223_o;
  wire [31:0] n224_o;
  wire n225_o;
  wire [31:0] n226_o;
  wire [31:0] n228_o;
  wire [31:0] n229_o;
  wire n233_o;
  wire n234_o;
  wire n235_o;
  wire n236_o;
  wire n240_o;
  wire [31:0] n241_o;
  wire n242_o;
  wire n243_o;
  wire [15:0] n245_o;
  wire [47:0] n246_o;
  wire [39:0] n247_o;
  wire [47:0] n249_o;
  wire [47:0] n250_o;
  wire n251_o;
  wire n252_o;
  wire [15:0] n253_o;
  wire n254_o;
  wire n255_o;
  wire [15:0] n256_o;
  wire [1:0] n257_o;
  wire n259_o;
  wire [7:0] n260_o;
  wire [7:0] n261_o;
  wire [15:0] n262_o;
  wire [1:0] n263_o;
  wire n265_o;
  wire [7:0] n266_o;
  wire [7:0] n267_o;
  wire [15:0] n268_o;
  wire [15:0] n269_o;
  wire [15:0] n270_o;
  wire [15:0] n271_o;
  wire [15:0] n272_o;
  wire [15:0] n273_o;
  wire n274_o;
  wire [7:0] n275_o;
  wire [7:0] n276_o;
  wire [15:0] n277_o;
  wire [15:0] n278_o;
  wire n291_o;
  wire n299_o;
  wire n302_o;
  wire n306_o;
  wire n316_o;
  wire n317_o;
  wire n318_o;
  wire n319_o;
  wire n320_o;
  wire [7:0] n325_o;
  wire [7:0] n326_o;
  wire [7:0] n327_o;
  wire [7:0] n328_o;
  wire [7:0] n329_o;
  wire [7:0] n330_o;
  wire [7:0] n331_o;
  wire [7:0] n332_o;
  wire [7:0] n333_o;
  wire [7:0] n334_o;
  wire [7:0] n335_o;
  wire [15:0] n336_o;
  wire [15:0] n337_o;
  wire [15:0] n338_o;
  wire [15:0] n339_o;
  wire [15:0] n340_o;
  wire [15:0] n341_o;
  wire [15:0] n342_o;
  wire [15:0] n343_o;
  wire [15:0] n344_o;
  wire [7:0] n345_o;
  wire [7:0] n346_o;
  wire [7:0] n347_o;
  wire [7:0] n348_o;
  wire [7:0] n349_o;
  wire [7:0] n350_o;
  wire [7:0] n351_o;
  wire [7:0] n352_o;
  wire [7:0] n353_o;
  wire n354_o;
  wire [15:0] n355_o;
  wire [15:0] n356_o;
  wire n357_o;
  wire n358_o;
  wire n359_o;
  wire n360_o;
  wire n361_o;
  wire n362_o;
  wire n364_o;
  wire n365_o;
  wire n368_o;
  wire n370_o;
  wire [1:0] n371_o;
  reg n374_o;
  reg n377_o;
  wire n380_o;
  wire n382_o;
  wire n384_o;
  wire n386_o;
  wire n388_o;
  wire n390_o;
  wire n392_o;
  wire n395_o;
  wire n398_o;
  wire n403_o;
  wire n404_o;
  wire [3:0] n405_o;
  wire n406_o;
  wire [2:0] n407_o;
  wire [3:0] n409_o;
  wire [2:0] n410_o;
  wire [3:0] n411_o;
  wire [3:0] n412_o;
  wire [2:0] n413_o;
  wire [3:0] n415_o;
  wire [2:0] n416_o;
  wire [3:0] n418_o;
  wire [2:0] n419_o;
  wire [3:0] n420_o;
  wire [2:0] n421_o;
  wire n423_o;
  wire n424_o;
  wire [2:0] n425_o;
  wire [3:0] n426_o;
  wire [2:0] n427_o;
  wire [3:0] n429_o;
  wire [3:0] n430_o;
  wire [3:0] n431_o;
  wire [3:0] n433_o;
  wire [3:0] n434_o;
  wire [3:0] n435_o;
  wire [3:0] n436_o;
  wire [3:0] n437_o;
  wire [3:0] n438_o;
  wire [3:0] n439_o;
  wire [3:0] n440_o;
  wire n444_o;
  wire n445_o;
  wire n446_o;
  wire [3:0] n448_o;
  wire [3:0] n449_o;
  wire [2:0] n450_o;
  wire [3:0] n452_o;
  wire [2:0] n453_o;
  wire [3:0] n455_o;
  wire [2:0] n456_o;
  wire [3:0] n458_o;
  wire [2:0] n459_o;
  wire [3:0] n461_o;
  wire [2:0] n462_o;
  wire [3:0] n464_o;
  wire [2:0] n465_o;
  wire [3:0] n466_o;
  wire n467_o;
  wire [2:0] n468_o;
  wire [3:0] n469_o;
  wire [3:0] n471_o;
  wire [3:0] n472_o;
  wire [3:0] n473_o;
  wire [3:0] n474_o;
  wire [3:0] n475_o;
  wire [3:0] n476_o;
  wire [3:0] n477_o;
  wire [3:0] n478_o;
  wire n482_o;
  wire n483_o;
  wire n484_o;
  wire n485_o;
  wire n486_o;
  wire n487_o;
  wire n488_o;
  wire n489_o;
  wire n490_o;
  wire [31:0] n491_o;
  wire [31:0] n492_o;
  wire [31:0] n494_o;
  wire [15:0] n498_o;
  wire n499_o;
  wire n500_o;
  wire n501_o;
  wire n502_o;
  wire n503_o;
  wire n504_o;
  wire n505_o;
  wire n506_o;
  wire n507_o;
  wire n508_o;
  wire n509_o;
  wire n510_o;
  wire n511_o;
  wire n512_o;
  wire n513_o;
  wire n514_o;
  wire [3:0] n515_o;
  wire [3:0] n516_o;
  wire [3:0] n517_o;
  wire [3:0] n518_o;
  wire [15:0] n519_o;
  wire n520_o;
  localparam [15:0] n521_o = 16'b1111111111111111;
  wire n522_o;
  wire n523_o;
  wire n524_o;
  wire n525_o;
  wire n526_o;
  wire n527_o;
  wire n528_o;
  wire n529_o;
  wire n530_o;
  wire n531_o;
  wire n532_o;
  wire [7:0] n533_o;
  wire n534_o;
  wire n535_o;
  wire n536_o;
  wire n537_o;
  wire n538_o;
  wire n539_o;
  wire n540_o;
  wire n541_o;
  wire [3:0] n542_o;
  wire [3:0] n543_o;
  wire [7:0] n544_o;
  wire n545_o;
  wire [2:0] n546_o;
  wire [2:0] n547_o;
  wire n549_o;
  wire n552_o;
  wire n555_o;
  wire n556_o;
  wire n557_o;
  wire n558_o;
  wire [15:0] n559_o;
  wire [15:0] n560_o;
  wire [15:0] n561_o;
  wire [15:0] n562_o;
  wire [15:0] n563_o;
  wire [31:0] n564_o;
  wire [15:0] n565_o;
  wire [15:0] n566_o;
  wire [15:0] n567_o;
  wire [15:0] n568_o;
  wire [15:0] n569_o;
  wire [31:0] n570_o;
  wire [31:0] n571_o;
  wire [31:0] n572_o;
  wire [15:0] n575_o;
  wire [15:0] n576_o;
  wire n577_o;
  wire n578_o;
  wire n579_o;
  wire n580_o;
  wire n581_o;
  wire n582_o;
  wire n583_o;
  wire n584_o;
  wire n585_o;
  wire n586_o;
  wire n587_o;
  wire n588_o;
  wire n589_o;
  wire n590_o;
  wire n591_o;
  wire n592_o;
  wire n593_o;
  wire n594_o;
  wire n595_o;
  wire n596_o;
  wire n597_o;
  wire n598_o;
  wire n599_o;
  wire n600_o;
  wire n601_o;
  wire [3:0] n602_o;
  wire [3:0] n603_o;
  wire [3:0] n604_o;
  wire [3:0] n605_o;
  wire [3:0] n606_o;
  wire [3:0] n607_o;
  wire [15:0] n608_o;
  wire [7:0] n609_o;
  wire [23:0] n610_o;
  wire [7:0] n611_o;
  wire [7:0] n612_o;
  wire [7:0] n613_o;
  wire [7:0] n614_o;
  wire [7:0] n615_o;
  wire [7:0] n616_o;
  wire [7:0] n617_o;
  wire [23:0] n618_o;
  wire [23:0] n619_o;
  wire [7:0] n620_o;
  wire [7:0] n621_o;
  wire [7:0] n622_o;
  wire [7:0] n623_o;
  wire [7:0] n624_o;
  wire [7:0] n625_o;
  wire [7:0] n626_o;
  wire n631_o;
  wire n633_o;
  wire n634_o;
  wire n635_o;
  wire n637_o;
  wire n639_o;
  wire n642_o;
  wire n644_o;
  wire n646_o;
  wire n647_o;
  wire n649_o;
  wire n650_o;
  wire n652_o;
  wire n654_o;
  wire n655_o;
  wire n656_o;
  wire n658_o;
  wire n660_o;
  wire n661_o;
  wire n663_o;
  wire n665_o;
  wire n667_o;
  wire n668_o;
  wire n670_o;
  wire n672_o;
  wire n673_o;
  wire n674_o;
  wire n675_o;
  wire n676_o;
  wire n677_o;
  wire n679_o;
  wire n680_o;
  wire n681_o;
  wire [31:0] n682_o;
  wire [31:0] n683_o;
  wire [31:0] n684_o;
  wire n685_o;
  wire n687_o;
  wire n689_o;
  wire n690_o;
  wire n692_o;
  wire n693_o;
  wire n694_o;
  wire n695_o;
  wire n696_o;
  wire n698_o;
  wire [11:0] n699_o;
  wire [15:0] n701_o;
  wire n702_o;
  wire [11:0] n703_o;
  wire [15:0] n705_o;
  wire n706_o;
  wire n707_o;
  wire n708_o;
  wire n709_o;
  wire [11:0] n710_o;
  wire [15:0] n712_o;
  wire n713_o;
  wire n714_o;
  wire n715_o;
  wire n716_o;
  wire [15:0] n717_o;
  wire n718_o;
  wire [15:0] n719_o;
  wire n720_o;
  wire n721_o;
  wire n722_o;
  wire n723_o;
  wire n724_o;
  wire n726_o;
  wire n727_o;
  wire n728_o;
  wire [23:0] n729_o;
  wire [23:0] n730_o;
  wire [23:0] n731_o;
  wire [7:0] n732_o;
  wire n733_o;
  wire [15:0] n734_o;
  wire [15:0] n735_o;
  wire [15:0] n736_o;
  wire [15:0] n737_o;
  wire [15:0] n738_o;
  wire [15:0] n739_o;
  wire [15:0] n740_o;
  wire [31:0] n741_o;
  wire [31:0] n742_o;
  wire [15:0] n743_o;
  wire [15:0] n744_o;
  wire [15:0] n745_o;
  wire [15:0] n746_o;
  wire [15:0] n747_o;
  wire [31:0] n748_o;
  wire [31:0] n749_o;
  wire [31:0] n750_o;
  wire [31:0] n751_o;
  wire [31:0] n752_o;
  wire [31:0] n753_o;
  wire [31:0] n754_o;
  wire [15:0] n755_o;
  wire [15:0] n756_o;
  wire [15:0] n757_o;
  wire [15:0] n758_o;
  wire [15:0] n759_o;
  wire n760_o;
  wire [31:0] n761_o;
  wire [31:0] n762_o;
  wire n763_o;
  wire n766_o;
  wire [31:0] n768_o;
  wire n769_o;
  wire n771_o;
  wire [31:0] n772_o;
  wire n773_o;
  wire n775_o;
  wire [31:0] n776_o;
  wire n777_o;
  wire n779_o;
  wire [31:0] n781_o;
  wire [31:0] n782_o;
  wire n783_o;
  wire n784_o;
  wire n785_o;
  wire n786_o;
  wire n787_o;
  wire n788_o;
  wire n789_o;
  wire [31:0] n790_o;
  wire [31:0] n791_o;
  wire n793_o;
  wire n795_o;
  wire n796_o;
  wire n798_o;
  wire n800_o;
  wire n801_o;
  wire n803_o;
  wire n816_o;
  wire [15:0] n817_o;
  wire n818_o;
  wire n819_o;
  wire n820_o;
  wire n821_o;
  wire n822_o;
  wire n823_o;
  wire n824_o;
  wire n825_o;
  wire n826_o;
  wire n827_o;
  wire n828_o;
  wire n829_o;
  wire n830_o;
  wire n831_o;
  wire n832_o;
  wire n833_o;
  wire [3:0] n834_o;
  wire [3:0] n835_o;
  wire [3:0] n836_o;
  wire [3:0] n837_o;
  wire [15:0] n838_o;
  wire [15:0] n839_o;
  wire [15:0] n840_o;
  wire [31:0] n841_o;
  wire n842_o;
  wire n844_o;
  wire n846_o;
  wire [1:0] n847_o;
  wire [15:0] n848_o;
  wire [31:0] n849_o;
  wire n851_o;
  wire [14:0] n852_o;
  wire [15:0] n853_o;
  wire [30:0] n854_o;
  wire [31:0] n856_o;
  wire n858_o;
  wire [13:0] n859_o;
  wire [15:0] n860_o;
  wire [29:0] n861_o;
  wire [31:0] n863_o;
  wire n865_o;
  wire [12:0] n866_o;
  wire [15:0] n867_o;
  wire [28:0] n868_o;
  wire [31:0] n870_o;
  wire n872_o;
  wire [3:0] n873_o;
  reg [31:0] n874_o;
  wire [31:0] n875_o;
  wire [9:0] n882_o;
  wire [9:0] n883_o;
  wire [9:0] n885_o;
  wire [9:0] n887_o;
  wire [9:0] n889_o;
  wire n890_o;
  wire [9:0] n892_o;
  wire [9:0] n894_o;
  wire [9:0] n896_o;
  wire [9:0] n898_o;
  wire [9:0] n900_o;
  wire [9:0] n902_o;
  wire [3:0] n903_o;
  wire [7:0] n905_o;
  wire [9:0] n907_o;
  wire [9:0] n908_o;
  wire n909_o;
  wire [9:0] n911_o;
  wire [9:0] n912_o;
  wire [31:0] n913_o;
  wire [31:0] n916_o;
  wire [31:0] n917_o;
  wire n919_o;
  wire n920_o;
  wire n921_o;
  wire [2:0] n922_o;
  wire n923_o;
  wire n924_o;
  wire n925_o;
  wire n926_o;
  wire n927_o;
  wire n928_o;
  wire n929_o;
  wire n930_o;
  wire [3:0] n931_o;
  wire [3:0] n932_o;
  wire [7:0] n933_o;
  wire n934_o;
  wire n935_o;
  wire n936_o;
  wire n937_o;
  wire n938_o;
  wire n939_o;
  wire n940_o;
  wire n941_o;
  wire n942_o;
  wire n943_o;
  wire n944_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n948_o;
  wire n949_o;
  wire [3:0] n950_o;
  wire [3:0] n951_o;
  wire [3:0] n952_o;
  wire [3:0] n953_o;
  wire [15:0] n954_o;
  wire n955_o;
  wire [31:0] n956_o;
  wire [7:0] n957_o;
  wire [7:0] n958_o;
  wire [7:0] n959_o;
  wire [23:0] n960_o;
  wire [23:0] n961_o;
  wire [23:0] n962_o;
  wire [31:0] n963_o;
  wire [31:0] n964_o;
  wire n965_o;
  wire n966_o;
  wire n969_o;
  wire n970_o;
  wire n971_o;
  wire n972_o;
  wire [4:0] n975_o;
  wire [4:0] n976_o;
  wire [3:0] n978_o;
  wire [4:0] n980_o;
  wire [4:0] n981_o;
  wire [4:0] n982_o;
  wire [4:0] n983_o;
  wire [4:0] n984_o;
  wire [26:0] n985_o;
  wire [26:0] n986_o;
  wire [26:0] n987_o;
  wire n989_o;
  wire n991_o;
  wire n992_o;
  wire n993_o;
  wire n994_o;
  wire n996_o;
  wire n997_o;
  wire n998_o;
  wire n999_o;
  wire n1000_o;
  wire n1001_o;
  wire n1002_o;
  wire n1004_o;
  wire n1005_o;
  wire n1006_o;
  wire n1008_o;
  wire n1009_o;
  wire n1010_o;
  wire n1011_o;
  wire n1012_o;
  wire n1015_o;
  wire [31:0] n1016_o;
  wire n1018_o;
  wire [31:0] n1019_o;
  wire [31:0] n1021_o;
  wire n1023_o;
  wire [31:0] n1024_o;
  wire [31:0] n1026_o;
  wire n1028_o;
  wire [31:0] n1029_o;
  wire [31:0] n1031_o;
  wire n1033_o;
  wire [31:0] n1034_o;
  wire [31:0] n1036_o;
  wire n1038_o;
  wire [31:0] n1039_o;
  wire [31:0] n1041_o;
  wire n1043_o;
  wire [31:0] n1044_o;
  wire [31:0] n1046_o;
  wire n1048_o;
  wire [31:0] n1049_o;
  wire [31:0] n1051_o;
  wire n1054_o;
  wire n1056_o;
  wire n1057_o;
  wire n1058_o;
  wire n1059_o;
  wire n1060_o;
  wire n1062_o;
  wire n1063_o;
  wire [31:0] n1072_o;
  wire [31:0] n1073_o;
  wire [31:0] n1074_o;
  wire n1075_o;
  wire [31:0] n1077_o;
  wire [31:0] n1081_o;
  localparam [2:0] n1082_o = 3'b000;
  wire n1083_o;
  wire n1084_o;
  wire n1085_o;
  wire n1086_o;
  wire n1087_o;
  wire [3:0] n1088_o;
  wire n1089_o;
  wire n1090_o;
  wire n1091_o;
  wire n1092_o;
  wire n1093_o;
  wire n1094_o;
  wire n1095_o;
  wire n1096_o;
  wire [3:0] n1097_o;
  wire [3:0] n1098_o;
  wire [7:0] n1099_o;
  wire n1100_o;
  wire n1101_o;
  wire n1102_o;
  wire n1103_o;
  wire n1104_o;
  wire n1105_o;
  wire n1106_o;
  wire n1107_o;
  wire n1108_o;
  wire n1109_o;
  wire n1110_o;
  wire n1111_o;
  wire n1112_o;
  wire n1113_o;
  wire n1114_o;
  wire n1115_o;
  wire [3:0] n1116_o;
  wire [3:0] n1117_o;
  wire [3:0] n1118_o;
  wire [3:0] n1119_o;
  wire [15:0] n1120_o;
  localparam [1:0] n1121_o = 2'b11;
  wire n1124_o;
  wire n1125_o;
  wire n1129_o;
  wire n1130_o;
  wire n1131_o;
  wire n1132_o;
  wire n1133_o;
  wire n1134_o;
  wire n1135_o;
  wire n1136_o;
  wire n1137_o;
  wire n1138_o;
  wire n1139_o;
  wire n1140_o;
  wire n1141_o;
  wire n1142_o;
  wire n1143_o;
  wire n1144_o;
  wire n1146_o;
  wire n1148_o;
  wire n1150_o;
  wire n1151_o;
  wire n1152_o;
  wire n1153_o;
  wire [2:0] n1154_o;
  wire n1155_o;
  wire n1156_o;
  wire [1:0] n1157_o;
  wire n1158_o;
  wire n1159_o;
  wire n1160_o;
  wire [1:0] n1161_o;
  wire [1:0] n1162_o;
  wire [7:0] n1166_o;
  wire [7:0] n1167_o;
  wire [7:0] n1168_o;
  wire [23:0] n1169_o;
  wire [23:0] n1170_o;
  wire [23:0] n1171_o;
  wire [31:0] n1172_o;
  wire [31:0] n1173_o;
  wire [31:0] n1174_o;
  wire [31:0] n1175_o;
  wire n1177_o;
  wire n1179_o;
  wire n1180_o;
  wire n1181_o;
  wire n1182_o;
  wire n1183_o;
  wire n1185_o;
  wire n1186_o;
  wire n1187_o;
  wire n1189_o;
  wire n1190_o;
  wire n1191_o;
  wire n1192_o;
  wire n1193_o;
  wire [2:0] n1194_o;
  wire n1195_o;
  wire n1197_o;
  wire n1198_o;
  wire n1199_o;
  wire n1200_o;
  wire n1201_o;
  wire n1204_o;
  wire n1206_o;
  wire n1209_o;
  wire n1211_o;
  wire n1215_o;
  wire n1218_o;
  wire n1221_o;
  wire n1223_o;
  wire n1224_o;
  wire n1225_o;
  wire n1226_o;
  wire n1227_o;
  wire n1229_o;
  wire n1230_o;
  wire n1231_o;
  wire n1232_o;
  wire n1233_o;
  wire n1236_o;
  wire [2:0] n1238_o;
  wire [3:0] n1240_o;
  wire [5:0] n1242_o;
  wire [1:0] n1243_o;
  wire [1:0] n1244_o;
  wire [3:0] n1245_o;
  wire n1246_o;
  wire n1247_o;
  wire n1249_o;
  wire n1250_o;
  wire n1251_o;
  wire n1252_o;
  wire [31:0] n1253_o;
  wire [31:0] n1254_o;
  wire [31:0] n1255_o;
  wire [31:0] n1256_o;
  wire [5:0] n1257_o;
  wire [3:0] n1258_o;
  wire n1259_o;
  wire n1260_o;
  wire n1262_o;
  wire n1263_o;
  wire n1264_o;
  wire n1265_o;
  wire [7:0] n1267_o;
  wire n1270_o;
  wire n1273_o;
  wire [2:0] n1274_o;
  wire [7:0] n1275_o;
  wire n1277_o;
  wire n1281_o;
  wire n1284_o;
  wire [2:0] n1286_o;
  wire [7:0] n1287_o;
  wire n1288_o;
  wire n1289_o;
  wire n1290_o;
  wire n1292_o;
  wire [2:0] n1293_o;
  wire [7:0] n1294_o;
  wire n1296_o;
  wire n1297_o;
  wire n1298_o;
  wire [7:0] n1299_o;
  wire [7:0] n1300_o;
  wire n1302_o;
  wire [15:0] n1303_o;
  wire [31:0] n1304_o;
  wire [15:0] n1305_o;
  wire [7:0] n1306_o;
  wire n1308_o;
  wire [7:0] n1309_o;
  wire n1311_o;
  wire n1312_o;
  wire n1313_o;
  wire n1315_o;
  wire n1317_o;
  wire n1319_o;
  wire n1321_o;
  wire n1323_o;
  wire n1324_o;
  wire [31:0] n1325_o;
  wire [31:0] n1326_o;
  wire [31:0] n1328_o;
  wire [5:0] n1329_o;
  wire [5:0] n1330_o;
  wire [31:0] n1331_o;
  wire [5:0] n1332_o;
  wire n1333_o;
  wire n1334_o;
  wire n1335_o;
  wire n1336_o;
  wire n1337_o;
  wire n1338_o;
  wire n1339_o;
  wire n1340_o;
  wire n1341_o;
  wire n1342_o;
  wire n1343_o;
  wire [1:0] n1345_o;
  wire [1:0] n1346_o;
  wire n1348_o;
  wire n1350_o;
  wire n1351_o;
  wire n1352_o;
  wire n1353_o;
  wire n1355_o;
  wire n1357_o;
  wire n1359_o;
  wire n1360_o;
  wire n1361_o;
  wire n1362_o;
  wire n1364_o;
  wire n1365_o;
  wire n1367_o;
  wire n1368_o;
  wire n1369_o;
  wire n1370_o;
  wire n1371_o;
  wire n1372_o;
  wire n1373_o;
  wire n1374_o;
  wire n1377_o;
  wire n1378_o;
  wire n1379_o;
  wire n1381_o;
  wire n1382_o;
  wire n1383_o;
  wire n1384_o;
  wire n1387_o;
  wire [5:0] n1390_o;
  wire [5:0] n1393_o;
  wire n1395_o;
  wire [5:0] n1397_o;
  wire [5:0] n1399_o;
  wire n1401_o;
  wire [5:0] n1402_o;
  wire [5:0] n1403_o;
  wire n1404_o;
  wire [5:0] n1406_o;
  wire [5:0] n1408_o;
  wire n1409_o;
  wire [1:0] n1410_o;
  wire [1:0] n1412_o;
  wire n1414_o;
  wire [5:0] n1415_o;
  wire [5:0] n1416_o;
  wire n1417_o;
  wire [1:0] n1418_o;
  wire [1:0] n1420_o;
  wire n1422_o;
  wire [5:0] n1424_o;
  wire [5:0] n1425_o;
  wire n1426_o;
  wire n1427_o;
  wire n1429_o;
  wire [1:0] n1430_o;
  wire n1431_o;
  wire n1432_o;
  wire n1434_o;
  wire n1435_o;
  wire [5:0] n1436_o;
  wire n1437_o;
  wire n1438_o;
  wire n1439_o;
  wire n1440_o;
  wire n1442_o;
  wire n1444_o;
  wire n1445_o;
  wire [15:0] n1446_o;
  wire [15:0] n1447_o;
  wire [15:0] n1448_o;
  wire n1449_o;
  wire n1450_o;
  wire n1452_o;
  wire [15:0] n1453_o;
  wire [15:0] n1454_o;
  wire [31:0] n1455_o;
  wire n1456_o;
  wire n1457_o;
  wire n1459_o;
  wire [15:0] n1461_o;
  wire n1463_o;
  wire [15:0] n1464_o;
  wire [31:0] n1465_o;
  wire n1467_o;
  wire n1468_o;
  wire [7:0] n1469_o;
  wire [1:0] n1470_o;
  wire [1:0] n1471_o;
  wire [1:0] n1472_o;
  wire [1:0] n1473_o;
  wire n1474_o;
  wire [15:0] n1475_o;
  wire [15:0] n1476_o;
  wire n1477_o;
  wire n1478_o;
  wire n1479_o;
  wire n1480_o;
  wire n1481_o;
  wire n1482_o;
  wire n1483_o;
  wire n1484_o;
  wire n1485_o;
  wire n1486_o;
  wire n1487_o;
  wire n1488_o;
  wire n1489_o;
  wire n1490_o;
  wire n1491_o;
  wire n1492_o;
  wire n1493_o;
  wire n1494_o;
  wire n1495_o;
  wire n1496_o;
  wire [7:0] n1497_o;
  wire n1498_o;
  wire n1499_o;
  wire [5:0] n1500_o;
  wire [3:0] n1502_o;
  wire [5:0] n1503_o;
  wire n1504_o;
  wire n1505_o;
  wire n1506_o;
  wire n1507_o;
  wire n1508_o;
  wire [1:0] n1509_o;
  wire [1:0] n1510_o;
  wire [31:0] n1512_o;
  wire [1:0] n1514_o;
  wire [1:0] n1515_o;
  wire n1517_o;
  wire [15:0] n1519_o;
  wire [15:0] n1520_o;
  wire [31:0] n1521_o;
  wire [31:0] n1522_o;
  wire [15:0] n1524_o;
  wire n1525_o;
  wire n1527_o;
  wire [15:0] n1528_o;
  wire n1530_o;
  wire n1532_o;
  wire n1534_o;
  wire n1536_o;
  wire n1538_o;
  wire [1:0] n1539_o;
  wire [5:0] n1541_o;
  wire n1543_o;
  wire n1545_o;
  wire n1547_o;
  wire [7:0] n1548_o;
  wire n1550_o;
  wire n1552_o;
  wire [2:0] n1553_o;
  wire [7:0] n1554_o;
  wire n1556_o;
  wire n1558_o;
  wire [5:0] n1560_o;
  wire [3:0] n1561_o;
  wire [5:0] n1562_o;
  wire n1563_o;
  wire [5:0] n1564_o;
  wire [5:0] n1565_o;
  wire [31:0] n1566_o;
  wire [5:0] n1567_o;
  wire n1608_o;
  wire n1609_o;
  wire n1610_o;
  wire n1611_o;
  wire n1612_o;
  wire n1614_o;
  wire n1615_o;
  wire n1617_o;
  wire n1618_o;
  wire n1619_o;
  wire n1620_o;
  wire n1623_o;
  wire n1624_o;
  wire n1625_o;
  wire [1:0] n1626_o;
  wire n1627_o;
  wire n1628_o;
  wire n1629_o;
  wire [35:0] n1630_o;
  wire [47:0] n1631_o;
  wire [88:0] n1632_o;
  wire n1633_o;
  wire n1634_o;
  wire n1635_o;
  wire n1636_o;
  wire n1637_o;
  wire [84:0] n1639_o;
  wire n1640_o;
  wire n1641_o;
  wire n1642_o;
  wire n1643_o;
  wire n1644_o;
  wire [1:0] n1645_o;
  wire n1647_o;
  wire [88:0] n1649_o;
  wire [88:0] n1650_o;
  wire n1652_o;
  wire n1653_o;
  wire [16:0] n1654_o;
  wire [16:0] n1655_o;
  wire [16:0] n1656_o;
  wire [70:0] n1657_o;
  wire [70:0] n1658_o;
  wire [70:0] n1659_o;
  wire [88:0] n1661_o;
  wire n1669_o;
  wire [4:0] n1670_o;
  wire [5:0] n1672_o;
  wire [4:0] n1673_o;
  wire [5:0] n1675_o;
  wire n1677_o;
  wire [4:0] n1678_o;
  localparam [31:0] n1679_o = 32'b00000000000000000000000000000000;
  wire [26:0] n1680_o;
  wire [31:0] n1681_o;
  wire [31:0] n1682_o;
  wire n1684_o;
  wire [4:0] n1685_o;
  wire [4:0] n1687_o;
  wire [4:0] n1688_o;
  wire [4:0] n1690_o;
  wire [4:0] n1691_o;
  wire [5:0] n1692_o;
  wire n1693_o;
  wire n1694_o;
  wire [2:0] n1695_o;
  wire n1697_o;
  wire [5:0] n1699_o;
  wire [4:0] n1702_o;
  wire [4:0] n1703_o;
  wire [4:0] n1704_o;
  wire [1:0] n1705_o;
  wire n1707_o;
  wire [2:0] n1708_o;
  wire n1710_o;
  wire [5:0] n1712_o;
  wire [5:0] n1714_o;
  wire [4:0] n1717_o;
  wire [4:0] n1718_o;
  wire [4:0] n1719_o;
  wire [2:0] n1720_o;
  wire n1722_o;
  wire [2:0] n1723_o;
  wire [5:0] n1725_o;
  wire [5:0] n1727_o;
  wire [4:0] n1729_o;
  wire [2:0] n1730_o;
  wire [2:0] n1732_o;
  wire [5:0] n1734_o;
  wire [5:0] n1735_o;
  wire [5:0] n1736_o;
  wire [1:0] n1738_o;
  wire [1:0] n1739_o;
  wire [1:0] n1740_o;
  wire [1:0] n1741_o;
  wire n1742_o;
  wire n1743_o;
  wire n1744_o;
  wire [2:0] n1745_o;
  wire [2:0] n1746_o;
  wire [2:0] n1747_o;
  wire [5:0] n1748_o;
  wire [5:0] n1749_o;
  wire [2:0] n1750_o;
  wire n1752_o;
  wire n1754_o;
  wire n1756_o;
  wire n1758_o;
  wire [3:0] n1759_o;
  reg [5:0] n1765_o;
  wire n1767_o;
  wire [5:0] n1769_o;
  wire n1773_o;
  wire [7:0] n1774_o;
  wire [7:0] n1775_o;
  wire n1776_o;
  wire [7:0] n1777_o;
  wire [7:0] n1778_o;
  wire n1779_o;
  wire [7:0] n1780_o;
  wire [7:0] n1781_o;
  wire [7:0] n1782_o;
  wire [7:0] n1783_o;
  wire [7:0] n1784_o;
  wire [7:0] n1785_o;
  wire n1788_o;
  wire n1789_o;
  wire n1790_o;
  wire n1791_o;
  wire n1792_o;
  wire n1793_o;
  wire n1794_o;
  wire n1795_o;
  wire n1796_o;
  wire n1797_o;
  wire n1798_o;
  wire n1800_o;
  wire n1801_o;
  wire n1803_o;
  wire n1804_o;
  wire n1805_o;
  wire n1806_o;
  wire n1807_o;
  wire n1808_o;
  wire n1809_o;
  wire n1810_o;
  wire n1811_o;
  wire n1812_o;
  wire n1814_o;
  wire n1816_o;
  wire n1818_o;
  wire n1819_o;
  wire n1821_o;
  wire n1822_o;
  wire n1823_o;
  wire [4:0] n1825_o;
  wire n1826_o;
  wire [7:0] n1827_o;
  wire n1829_o;
  wire [2:0] n1830_o;
  wire [2:0] n1831_o;
  wire [2:0] n1832_o;
  wire [2:0] n1833_o;
  wire [4:0] n1834_o;
  wire [4:0] n1835_o;
  wire [4:0] n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1839_o;
  wire n1840_o;
  wire n1841_o;
  wire n1842_o;
  wire [7:0] n1843_o;
  wire n1846_o;
  wire n1847_o;
  wire n1848_o;
  wire n1851_o;
  wire n1852_o;
  wire n1853_o;
  wire n1854_o;
  wire n1855_o;
  wire n1856_o;
  wire n1857_o;
  wire n1858_o;
  wire n1865_o;
  wire n1866_o;
  wire n1867_o;
  wire n1868_o;
  wire n1869_o;
  wire n1870_o;
  wire [2:0] n1872_o;
  wire [2:0] n1873_o;
  wire [2:0] n1874_o;
  wire n1875_o;
  wire n1876_o;
  wire [7:0] n1877_o;
  wire [7:0] n1878_o;
  wire n1879_o;
  wire n1880_o;
  wire n1881_o;
  wire n1882_o;
  wire [7:0] n1884_o;
  wire n1886_o;
  wire n1888_o;
  wire n1890_o;
  wire [1:0] n1900_o;
  wire n1902_o;
  wire [5:0] n1904_o;
  wire [5:0] n1906_o;
  localparam [88:0] n1909_o = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [1:0] n1912_o;
  wire n1914_o;
  wire n1916_o;
  wire [1:0] n1917_o;
  reg [1:0] n1921_o;
  wire n1922_o;
  wire n1924_o;
  wire n1925_o;
  wire n1928_o;
  wire n1929_o;
  wire n1931_o;
  wire n1932_o;
  wire [1:0] n1935_o;
  wire n1938_o;
  wire [1:0] n1940_o;
  wire [6:0] n1943_o;
  wire n1945_o;
  wire n1946_o;
  wire n1947_o;
  wire n1948_o;
  wire n1949_o;
  wire n1950_o;
  wire n1951_o;
  wire [6:0] n1954_o;
  wire [6:0] n1956_o;
  wire n1957_o;
  wire n1959_o;
  wire n1960_o;
  wire n1961_o;
  wire n1963_o;
  wire [1:0] n1965_o;
  wire n1967_o;
  wire n1968_o;
  wire [6:0] n1971_o;
  wire n1973_o;
  wire n1974_o;
  wire n1975_o;
  wire n1976_o;
  wire n1977_o;
  wire [6:0] n1980_o;
  wire n1981_o;
  wire n1983_o;
  wire [1:0] n1985_o;
  wire n1986_o;
  wire [6:0] n1987_o;
  wire n1989_o;
  wire n1990_o;
  wire n1991_o;
  wire n1992_o;
  wire n1994_o;
  wire [1:0] n1996_o;
  wire n1997_o;
  wire n1998_o;
  wire n1999_o;
  wire n2000_o;
  wire n2002_o;
  wire n2003_o;
  wire [1:0] n2006_o;
  wire n2007_o;
  wire [6:0] n2009_o;
  wire n2010_o;
  wire n2015_o;
  wire [1:0] n2017_o;
  wire [1:0] n2018_o;
  wire [1:0] n2019_o;
  wire n2022_o;
  wire n2023_o;
  wire n2024_o;
  wire [1:0] n2026_o;
  wire n2027_o;
  wire n2028_o;
  wire n2029_o;
  wire n2031_o;
  wire n2032_o;
  wire n2035_o;
  wire n2036_o;
  wire n2037_o;
  wire [2:0] n2038_o;
  wire n2040_o;
  wire [2:0] n2042_o;
  wire n2044_o;
  wire n2046_o;
  wire n2047_o;
  wire n2048_o;
  wire n2049_o;
  wire n2051_o;
  wire n2052_o;
  wire [2:0] n2054_o;
  wire n2056_o;
  wire n2058_o;
  wire n2059_o;
  wire n2060_o;
  wire n2061_o;
  wire n2063_o;
  wire n2065_o;
  wire n2066_o;
  wire n2068_o;
  wire n2069_o;
  wire n2071_o;
  wire n2073_o;
  wire [2:0] n2074_o;
  wire n2076_o;
  wire n2079_o;
  wire n2082_o;
  wire n2085_o;
  wire n2087_o;
  wire n2089_o;
  wire n2091_o;
  wire [4:0] n2092_o;
  reg n2095_o;
  reg n2098_o;
  reg n2101_o;
  reg n2105_o;
  reg n2109_o;
  wire n2110_o;
  reg n2111_o;
  reg n2112_o;
  reg [6:0] n2117_o;
  wire n2119_o;
  wire [3:0] n2120_o;
  reg n2123_o;
  reg n2126_o;
  reg n2128_o;
  reg n2130_o;
  reg n2132_o;
  wire n2133_o;
  reg n2134_o;
  wire n2135_o;
  reg n2136_o;
  wire n2137_o;
  reg n2138_o;
  wire n2139_o;
  reg n2140_o;
  wire n2141_o;
  reg n2142_o;
  reg n2143_o;
  reg [6:0] n2146_o;
  wire n2148_o;
  wire n2151_o;
  wire n2154_o;
  wire n2157_o;
  wire n2160_o;
  wire [1:0] n2162_o;
  wire n2163_o;
  wire n2164_o;
  wire [1:0] n2165_o;
  wire [1:0] n2166_o;
  wire n2167_o;
  wire n2168_o;
  wire n2169_o;
  wire n2170_o;
  wire n2171_o;
  wire [1:0] n2177_o;
  wire [1:0] n2178_o;
  wire [10:0] n2179_o;
  wire [6:0] n2180_o;
  wire n2181_o;
  wire n2183_o;
  wire n2184_o;
  wire [3:0] n2185_o;
  wire n2186_o;
  wire [2:0] n2187_o;
  wire n2189_o;
  wire n2190_o;
  wire n2193_o;
  wire n2194_o;
  wire n2198_o;
  wire n2199_o;
  wire n2201_o;
  wire n2203_o;
  wire n2204_o;
  wire n2206_o;
  wire n2207_o;
  wire n2208_o;
  wire n2210_o;
  wire n2211_o;
  wire n2212_o;
  wire [6:0] n2214_o;
  wire n2217_o;
  wire n2218_o;
  wire [2:0] n2219_o;
  wire n2221_o;
  wire n2222_o;
  wire [2:0] n2223_o;
  wire n2225_o;
  wire [5:0] n2226_o;
  wire n2228_o;
  wire n2229_o;
  wire n2230_o;
  wire n2231_o;
  wire n2232_o;
  wire [6:0] n2233_o;
  wire n2235_o;
  wire [1:0] n2236_o;
  wire n2238_o;
  wire n2239_o;
  wire n2240_o;
  wire [1:0] n2241_o;
  wire n2243_o;
  wire [2:0] n2244_o;
  wire n2246_o;
  wire n2247_o;
  wire [1:0] n2248_o;
  wire n2250_o;
  wire n2251_o;
  wire n2252_o;
  wire [1:0] n2255_o;
  wire n2257_o;
  wire [1:0] n2258_o;
  wire n2260_o;
  wire n2263_o;
  wire n2266_o;
  wire n2268_o;
  wire [1:0] n2269_o;
  wire n2271_o;
  wire [1:0] n2274_o;
  wire n2275_o;
  wire n2276_o;
  wire n2279_o;
  wire n2280_o;
  wire n2281_o;
  wire n2282_o;
  wire [6:0] n2284_o;
  wire n2287_o;
  wire n2289_o;
  wire n2291_o;
  wire n2292_o;
  wire [1:0] n2293_o;
  wire n2295_o;
  wire n2298_o;
  wire n2301_o;
  wire n2303_o;
  wire n2305_o;
  wire n2307_o;
  wire n2309_o;
  wire n2311_o;
  wire n2313_o;
  wire n2314_o;
  wire [2:0] n2315_o;
  wire n2317_o;
  wire n2318_o;
  wire n2319_o;
  wire [1:0] n2320_o;
  wire n2322_o;
  wire [1:0] n2323_o;
  wire n2325_o;
  wire n2326_o;
  wire [2:0] n2327_o;
  wire n2329_o;
  wire [1:0] n2330_o;
  wire n2332_o;
  wire n2333_o;
  wire n2334_o;
  wire n2335_o;
  wire [5:0] n2336_o;
  wire n2338_o;
  wire n2339_o;
  wire n2340_o;
  wire [1:0] n2341_o;
  wire n2343_o;
  wire n2345_o;
  wire [1:0] n2346_o;
  reg [1:0] n2350_o;
  wire n2351_o;
  wire [5:0] n2352_o;
  wire n2354_o;
  wire n2355_o;
  wire n2357_o;
  wire n2358_o;
  wire [6:0] n2360_o;
  wire n2363_o;
  wire n2364_o;
  wire n2365_o;
  wire n2366_o;
  wire [6:0] n2368_o;
  wire n2370_o;
  wire n2371_o;
  wire [1:0] n2377_o;
  wire n2380_o;
  wire n2381_o;
  wire n2382_o;
  wire n2383_o;
  wire n2384_o;
  wire n2385_o;
  wire n2386_o;
  wire n2387_o;
  wire n2388_o;
  wire [6:0] n2390_o;
  wire [1:0] n2391_o;
  wire n2393_o;
  wire n2394_o;
  wire n2395_o;
  wire n2396_o;
  wire n2397_o;
  wire n2398_o;
  wire n2399_o;
  wire n2400_o;
  wire n2401_o;
  wire n2402_o;
  wire n2403_o;
  wire n2404_o;
  wire [6:0] n2405_o;
  wire [1:0] n2406_o;
  wire [1:0] n2407_o;
  wire n2409_o;
  wire n2412_o;
  wire n2415_o;
  wire n2416_o;
  wire n2417_o;
  wire n2418_o;
  wire n2419_o;
  wire n2420_o;
  wire n2421_o;
  wire n2422_o;
  wire n2423_o;
  wire n2424_o;
  wire n2425_o;
  wire n2426_o;
  wire n2427_o;
  wire [6:0] n2428_o;
  wire [1:0] n2429_o;
  wire n2431_o;
  wire [1:0] n2432_o;
  wire n2434_o;
  wire n2435_o;
  wire [2:0] n2436_o;
  wire n2438_o;
  wire n2439_o;
  wire [2:0] n2440_o;
  wire n2442_o;
  wire n2443_o;
  wire [3:0] n2444_o;
  wire n2446_o;
  wire n2447_o;
  wire [1:0] n2449_o;
  wire n2452_o;
  wire n2453_o;
  wire n2454_o;
  wire n2455_o;
  wire [6:0] n2457_o;
  wire n2458_o;
  wire n2461_o;
  wire n2462_o;
  wire n2463_o;
  wire n2464_o;
  wire n2466_o;
  wire n2467_o;
  wire n2470_o;
  wire n2473_o;
  wire [1:0] n2475_o;
  wire n2477_o;
  wire n2478_o;
  wire n2479_o;
  wire [6:0] n2481_o;
  wire [1:0] n2482_o;
  wire n2483_o;
  wire n2486_o;
  wire n2489_o;
  wire n2491_o;
  wire [1:0] n2492_o;
  wire n2494_o;
  wire [1:0] n2495_o;
  wire [1:0] n2496_o;
  wire n2498_o;
  wire n2500_o;
  wire n2502_o;
  wire [6:0] n2503_o;
  wire [1:0] n2504_o;
  wire [1:0] n2505_o;
  wire n2507_o;
  wire n2508_o;
  wire n2509_o;
  wire n2511_o;
  wire n2513_o;
  wire n2514_o;
  wire n2515_o;
  wire n2516_o;
  wire n2517_o;
  wire n2518_o;
  wire n2519_o;
  wire n2520_o;
  wire n2521_o;
  wire n2522_o;
  wire n2524_o;
  wire n2525_o;
  wire n2526_o;
  wire n2527_o;
  wire n2529_o;
  wire n2531_o;
  wire [6:0] n2532_o;
  wire [1:0] n2533_o;
  wire [1:0] n2534_o;
  wire n2536_o;
  wire n2538_o;
  wire n2540_o;
  wire n2542_o;
  wire [1:0] n2543_o;
  wire [1:0] n2544_o;
  wire n2546_o;
  wire n2547_o;
  wire n2548_o;
  wire [1:0] n2549_o;
  wire [1:0] n2550_o;
  wire [1:0] n2551_o;
  wire [1:0] n2552_o;
  wire n2553_o;
  wire n2554_o;
  wire n2555_o;
  wire n2556_o;
  wire n2558_o;
  wire n2560_o;
  wire [6:0] n2561_o;
  wire [2:0] n2562_o;
  wire n2564_o;
  wire n2565_o;
  wire [1:0] n2566_o;
  wire n2568_o;
  wire n2569_o;
  wire [1:0] n2570_o;
  wire n2572_o;
  wire n2573_o;
  wire [2:0] n2574_o;
  wire n2576_o;
  wire [1:0] n2577_o;
  wire n2579_o;
  wire n2580_o;
  wire n2581_o;
  wire n2584_o;
  wire n2587_o;
  wire n2589_o;
  wire n2591_o;
  wire [1:0] n2592_o;
  wire n2594_o;
  wire [2:0] n2595_o;
  wire n2597_o;
  wire n2598_o;
  wire [2:0] n2599_o;
  wire n2601_o;
  wire [2:0] n2602_o;
  wire n2604_o;
  wire [1:0] n2605_o;
  wire n2607_o;
  wire n2608_o;
  wire [2:0] n2609_o;
  wire n2611_o;
  wire n2612_o;
  wire n2613_o;
  wire n2614_o;
  wire n2615_o;
  wire n2619_o;
  wire n2622_o;
  wire n2624_o;
  wire n2626_o;
  wire n2628_o;
  wire n2630_o;
  wire [2:0] n2631_o;
  wire n2633_o;
  wire [2:0] n2634_o;
  wire n2636_o;
  wire [1:0] n2637_o;
  wire n2639_o;
  wire n2640_o;
  wire [2:0] n2641_o;
  wire n2643_o;
  wire n2644_o;
  wire n2645_o;
  wire n2646_o;
  wire n2647_o;
  wire n2650_o;
  wire n2652_o;
  wire n2654_o;
  wire n2655_o;
  wire n2656_o;
  wire n2658_o;
  wire [2:0] n2659_o;
  wire n2661_o;
  wire [2:0] n2662_o;
  wire n2664_o;
  wire n2665_o;
  wire [2:0] n2666_o;
  wire n2668_o;
  wire [1:0] n2669_o;
  wire n2671_o;
  wire n2672_o;
  wire n2675_o;
  wire n2677_o;
  wire n2679_o;
  wire n2680_o;
  wire n2681_o;
  wire n2683_o;
  wire [2:0] n2684_o;
  wire n2686_o;
  wire [2:0] n2687_o;
  wire n2689_o;
  wire [1:0] n2690_o;
  wire n2692_o;
  wire n2693_o;
  wire [2:0] n2694_o;
  wire n2696_o;
  wire n2697_o;
  wire n2698_o;
  wire n2699_o;
  wire n2700_o;
  wire n2703_o;
  wire n2705_o;
  wire n2707_o;
  wire n2708_o;
  wire n2709_o;
  wire n2711_o;
  wire [2:0] n2712_o;
  wire n2714_o;
  wire [2:0] n2715_o;
  wire n2717_o;
  wire n2718_o;
  wire n2719_o;
  wire n2720_o;
  wire n2723_o;
  wire n2725_o;
  wire n2727_o;
  wire n2728_o;
  wire n2729_o;
  wire n2731_o;
  wire n2732_o;
  wire n2733_o;
  wire n2734_o;
  wire n2735_o;
  wire n2736_o;
  wire n2737_o;
  wire n2738_o;
  wire n2739_o;
  wire n2740_o;
  wire n2741_o;
  wire n2742_o;
  wire [5:0] n2743_o;
  wire n2745_o;
  wire n2746_o;
  wire n2747_o;
  wire n2748_o;
  wire n2749_o;
  wire n2750_o;
  wire n2751_o;
  wire n2752_o;
  wire n2753_o;
  wire n2754_o;
  wire n2755_o;
  wire n2756_o;
  wire n2758_o;
  wire n2760_o;
  wire n2761_o;
  wire n2763_o;
  wire n2764_o;
  wire n2765_o;
  wire [1:0] n2767_o;
  wire [2:0] n2768_o;
  wire [1:0] n2769_o;
  wire [2:0] n2770_o;
  wire [2:0] n2771_o;
  wire [1:0] n2772_o;
  wire [1:0] n2773_o;
  wire [6:0] n2775_o;
  wire [1:0] n2776_o;
  wire n2779_o;
  wire n2781_o;
  wire [2:0] n2782_o;
  wire [2:0] n2783_o;
  wire n2784_o;
  wire n2785_o;
  wire [1:0] n2786_o;
  wire [1:0] n2787_o;
  wire [6:0] n2788_o;
  wire n2789_o;
  wire n2790_o;
  wire [5:0] n2791_o;
  wire n2793_o;
  wire n2794_o;
  wire n2795_o;
  wire n2796_o;
  wire n2797_o;
  wire n2798_o;
  wire n2799_o;
  wire n2800_o;
  wire n2801_o;
  wire n2805_o;
  wire n2807_o;
  wire n2809_o;
  wire n2810_o;
  wire n2811_o;
  wire n2812_o;
  wire n2813_o;
  wire n2814_o;
  wire [6:0] n2816_o;
  wire [1:0] n2817_o;
  wire n2819_o;
  wire n2822_o;
  wire [2:0] n2823_o;
  wire n2825_o;
  wire [1:0] n2826_o;
  wire n2828_o;
  wire n2831_o;
  wire n2834_o;
  wire n2836_o;
  wire [1:0] n2837_o;
  wire n2839_o;
  wire n2841_o;
  wire n2842_o;
  wire n2844_o;
  wire n2845_o;
  wire n2847_o;
  wire n2849_o;
  wire n2851_o;
  wire n2853_o;
  wire n2855_o;
  wire n2856_o;
  wire n2858_o;
  wire n2860_o;
  wire n2861_o;
  wire [1:0] n2862_o;
  wire n2864_o;
  wire n2865_o;
  wire n2866_o;
  wire n2868_o;
  wire n2869_o;
  wire [2:0] n2870_o;
  wire [2:0] n2871_o;
  wire n2872_o;
  wire n2873_o;
  wire n2874_o;
  wire n2875_o;
  wire [1:0] n2876_o;
  wire [1:0] n2877_o;
  wire n2878_o;
  wire n2879_o;
  wire n2880_o;
  wire n2881_o;
  wire n2882_o;
  wire n2884_o;
  wire n2886_o;
  wire [6:0] n2887_o;
  wire n2888_o;
  wire n2890_o;
  wire n2891_o;
  wire n2893_o;
  wire n2895_o;
  wire n2897_o;
  wire n2899_o;
  wire n2900_o;
  wire n2901_o;
  wire n2903_o;
  wire n2905_o;
  wire n2906_o;
  wire n2907_o;
  wire n2908_o;
  wire n2909_o;
  wire n2910_o;
  wire n2912_o;
  wire n2914_o;
  wire [6:0] n2915_o;
  wire n2916_o;
  wire n2918_o;
  wire n2919_o;
  wire n2921_o;
  wire n2923_o;
  wire n2925_o;
  wire n2927_o;
  wire n2929_o;
  wire n2931_o;
  wire n2933_o;
  wire n2935_o;
  wire n2937_o;
  wire n2938_o;
  wire [3:0] n2939_o;
  wire n2941_o;
  wire [3:0] n2943_o;
  wire n2945_o;
  wire n2947_o;
  wire n2948_o;
  wire [1:0] n2949_o;
  wire n2951_o;
  wire n2952_o;
  wire n2953_o;
  wire n2954_o;
  wire n2956_o;
  wire [2:0] n2957_o;
  wire [2:0] n2958_o;
  wire n2959_o;
  wire n2960_o;
  wire n2961_o;
  wire n2962_o;
  wire [1:0] n2963_o;
  wire [1:0] n2964_o;
  wire n2965_o;
  wire n2966_o;
  wire n2967_o;
  wire n2968_o;
  wire n2969_o;
  wire n2971_o;
  wire [3:0] n2973_o;
  wire n2975_o;
  wire n2977_o;
  wire [6:0] n2978_o;
  wire n2979_o;
  wire [1:0] n2980_o;
  wire n2982_o;
  wire n2984_o;
  wire n2985_o;
  wire n2986_o;
  wire n2988_o;
  wire n2989_o;
  wire n2991_o;
  wire [2:0] n2992_o;
  wire [2:0] n2993_o;
  wire n2995_o;
  wire n2997_o;
  wire n2998_o;
  wire n2999_o;
  wire n3000_o;
  wire n3001_o;
  wire n3002_o;
  wire n3003_o;
  wire n3004_o;
  wire [1:0] n3005_o;
  wire [1:0] n3006_o;
  wire n3007_o;
  wire n3008_o;
  wire n3009_o;
  wire n3010_o;
  wire n3011_o;
  wire n3012_o;
  wire n3013_o;
  wire n3015_o;
  wire n3017_o;
  wire n3019_o;
  wire n3021_o;
  wire [3:0] n3023_o;
  wire n3025_o;
  wire n3027_o;
  wire [6:0] n3028_o;
  wire [1:0] n3029_o;
  wire [1:0] n3030_o;
  wire n3031_o;
  wire n3033_o;
  wire n3034_o;
  wire n3035_o;
  wire n3037_o;
  wire n3038_o;
  wire n3040_o;
  wire n3042_o;
  wire [1:0] n3043_o;
  wire [1:0] n3044_o;
  wire [2:0] n3045_o;
  wire [2:0] n3046_o;
  wire n3047_o;
  wire n3048_o;
  wire n3049_o;
  wire n3050_o;
  wire n3051_o;
  wire n3052_o;
  wire n3053_o;
  wire n3054_o;
  wire n3055_o;
  wire n3056_o;
  wire n3057_o;
  wire [1:0] n3058_o;
  wire [1:0] n3059_o;
  wire [1:0] n3060_o;
  wire [1:0] n3061_o;
  wire n3062_o;
  wire n3063_o;
  wire n3064_o;
  wire n3065_o;
  wire n3066_o;
  wire n3067_o;
  wire n3068_o;
  wire n3069_o;
  wire n3071_o;
  wire [3:0] n3073_o;
  wire n3075_o;
  wire n3076_o;
  wire n3077_o;
  wire [6:0] n3078_o;
  wire [1:0] n3080_o;
  wire [1:0] n3081_o;
  wire n3083_o;
  wire n3085_o;
  wire n3087_o;
  wire n3088_o;
  wire n3090_o;
  wire n3092_o;
  wire n3094_o;
  wire n3096_o;
  wire n3098_o;
  wire [1:0] n3099_o;
  wire [1:0] n3100_o;
  wire [2:0] n3101_o;
  wire [2:0] n3102_o;
  wire n3103_o;
  wire n3104_o;
  wire n3105_o;
  wire n3106_o;
  wire n3107_o;
  wire n3108_o;
  wire [1:0] n3109_o;
  wire [1:0] n3110_o;
  wire n3111_o;
  wire n3112_o;
  wire n3113_o;
  wire n3114_o;
  wire [1:0] n3115_o;
  wire [1:0] n3116_o;
  wire [1:0] n3117_o;
  wire [1:0] n3118_o;
  wire n3119_o;
  wire n3120_o;
  wire n3121_o;
  wire n3122_o;
  wire n3123_o;
  wire n3124_o;
  wire n3125_o;
  wire n3126_o;
  wire n3127_o;
  wire n3129_o;
  wire n3131_o;
  wire [3:0] n3133_o;
  wire n3135_o;
  wire n3137_o;
  wire n3138_o;
  wire [6:0] n3139_o;
  wire n3141_o;
  wire [1:0] n3142_o;
  wire n3144_o;
  wire [2:0] n3145_o;
  wire n3147_o;
  wire n3148_o;
  wire [3:0] n3149_o;
  wire n3151_o;
  wire [1:0] n3152_o;
  wire n3154_o;
  wire n3155_o;
  wire n3156_o;
  wire n3157_o;
  wire [2:0] n3158_o;
  wire n3160_o;
  wire [2:0] n3161_o;
  wire n3163_o;
  wire n3164_o;
  wire n3165_o;
  wire n3166_o;
  wire [2:0] n3168_o;
  wire n3170_o;
  wire n3172_o;
  wire n3173_o;
  wire [1:0] n3174_o;
  wire n3176_o;
  wire [1:0] n3177_o;
  wire n3179_o;
  wire n3182_o;
  wire n3184_o;
  wire [1:0] n3185_o;
  wire n3187_o;
  wire n3189_o;
  wire [1:0] n3190_o;
  reg [1:0] n3194_o;
  wire n3195_o;
  wire n3198_o;
  wire [1:0] n3199_o;
  wire n3201_o;
  wire n3202_o;
  wire [2:0] n3203_o;
  wire n3205_o;
  wire n3208_o;
  wire n3210_o;
  wire n3213_o;
  wire n3215_o;
  wire [1:0] n3216_o;
  wire n3218_o;
  wire n3219_o;
  wire n3220_o;
  wire n3221_o;
  wire [2:0] n3222_o;
  wire n3225_o;
  wire n3227_o;
  wire n3228_o;
  wire n3229_o;
  wire [2:0] n3231_o;
  wire n3233_o;
  wire n3235_o;
  wire n3236_o;
  wire n3237_o;
  wire n3238_o;
  wire n3239_o;
  wire n3240_o;
  wire n3241_o;
  wire [2:0] n3243_o;
  wire n3245_o;
  wire n3247_o;
  wire n3248_o;
  wire n3249_o;
  wire n3250_o;
  wire n3251_o;
  wire n3252_o;
  wire n3253_o;
  wire n3255_o;
  wire n3256_o;
  wire n3258_o;
  wire n3260_o;
  wire n3261_o;
  wire n3263_o;
  wire n3264_o;
  wire n3266_o;
  wire n3268_o;
  wire [2:0] n3269_o;
  wire n3271_o;
  wire n3274_o;
  wire [1:0] n3275_o;
  reg n3276_o;
  reg [6:0] n3279_o;
  wire n3281_o;
  wire [4:0] n3282_o;
  reg [1:0] n3284_o;
  reg n3286_o;
  wire n3287_o;
  reg n3288_o;
  wire n3289_o;
  wire n3290_o;
  wire n3291_o;
  reg n3292_o;
  wire n3293_o;
  wire n3294_o;
  wire n3295_o;
  reg n3296_o;
  reg n3297_o;
  reg n3298_o;
  reg n3299_o;
  reg [6:0] n3303_o;
  wire [1:0] n3304_o;
  wire n3305_o;
  wire [1:0] n3306_o;
  wire n3307_o;
  wire n3308_o;
  wire [1:0] n3309_o;
  wire n3310_o;
  wire n3311_o;
  wire n3312_o;
  wire [6:0] n3313_o;
  wire [1:0] n3314_o;
  wire n3315_o;
  wire n3316_o;
  wire n3318_o;
  wire n3321_o;
  wire n3323_o;
  wire n3325_o;
  wire n3328_o;
  wire n3331_o;
  wire n3334_o;
  wire [1:0] n3335_o;
  wire n3337_o;
  wire n3338_o;
  wire n3339_o;
  wire [1:0] n3340_o;
  wire [1:0] n3341_o;
  wire n3342_o;
  wire n3344_o;
  wire n3346_o;
  wire n3347_o;
  wire n3349_o;
  wire n3351_o;
  wire n3352_o;
  wire n3354_o;
  wire n3355_o;
  wire n3356_o;
  wire n3357_o;
  wire [2:0] n3358_o;
  wire n3360_o;
  wire [2:0] n3361_o;
  wire n3363_o;
  wire n3364_o;
  wire n3365_o;
  wire n3366_o;
  wire n3367_o;
  wire n3374_o;
  wire n3377_o;
  wire n3380_o;
  wire n3382_o;
  wire n3384_o;
  wire n3386_o;
  wire n3388_o;
  wire n3389_o;
  wire n3390_o;
  wire [1:0] n3391_o;
  wire n3393_o;
  wire n3394_o;
  wire n3395_o;
  wire [2:0] n3396_o;
  wire n3398_o;
  wire n3399_o;
  wire [3:0] n3400_o;
  wire n3402_o;
  wire n3403_o;
  wire [2:0] n3407_o;
  wire n3409_o;
  wire n3412_o;
  wire n3415_o;
  wire n3418_o;
  wire n3419_o;
  wire [1:0] n3421_o;
  wire n3423_o;
  wire n3425_o;
  wire n3427_o;
  wire n3428_o;
  wire n3431_o;
  wire n3434_o;
  wire n3437_o;
  wire n3439_o;
  wire n3441_o;
  wire n3442_o;
  wire n3445_o;
  wire n3448_o;
  wire n3450_o;
  wire n3451_o;
  wire n3452_o;
  wire n3454_o;
  wire n3456_o;
  wire [1:0] n3457_o;
  wire n3459_o;
  wire n3461_o;
  wire n3462_o;
  wire n3464_o;
  wire n3466_o;
  wire n3467_o;
  wire n3468_o;
  wire n3469_o;
  wire n3471_o;
  wire n3472_o;
  wire n3473_o;
  wire n3474_o;
  wire n3476_o;
  wire n3477_o;
  wire n3479_o;
  wire [2:0] n3480_o;
  wire n3482_o;
  wire [3:0] n3483_o;
  wire n3485_o;
  wire [1:0] n3486_o;
  wire n3488_o;
  wire n3489_o;
  wire n3490_o;
  wire n3491_o;
  wire n3493_o;
  wire n3494_o;
  wire n3495_o;
  wire n3496_o;
  wire n3497_o;
  wire n3498_o;
  wire n3499_o;
  wire n3500_o;
  wire n3503_o;
  wire n3504_o;
  wire n3506_o;
  wire n3507_o;
  wire n3508_o;
  wire n3509_o;
  wire n3510_o;
  wire n3511_o;
  wire n3512_o;
  wire n3513_o;
  wire n3516_o;
  wire [1:0] n3518_o;
  wire n3521_o;
  wire n3523_o;
  wire n3524_o;
  wire n3525_o;
  wire [1:0] n3527_o;
  wire n3529_o;
  wire n3530_o;
  wire n3531_o;
  wire n3532_o;
  wire n3533_o;
  wire n3534_o;
  wire [1:0] n3535_o;
  wire n3537_o;
  wire n3538_o;
  wire n3539_o;
  wire n3540_o;
  wire n3541_o;
  wire n3543_o;
  wire n3544_o;
  wire n3547_o;
  wire n3551_o;
  wire n3554_o;
  wire n3556_o;
  wire n3558_o;
  wire n3561_o;
  wire n3562_o;
  wire n3563_o;
  wire n3565_o;
  wire [1:0] n3566_o;
  wire n3568_o;
  wire n3570_o;
  wire n3572_o;
  wire n3574_o;
  wire n3576_o;
  wire n3577_o;
  wire n3578_o;
  wire n3580_o;
  wire n3582_o;
  wire [1:0] n3583_o;
  wire [1:0] n3584_o;
  wire n3586_o;
  wire n3588_o;
  wire n3589_o;
  wire n3591_o;
  wire n3592_o;
  wire n3593_o;
  wire n3594_o;
  wire n3595_o;
  wire n3596_o;
  wire n3597_o;
  wire n3598_o;
  wire n3599_o;
  wire n3600_o;
  wire n3601_o;
  wire n3602_o;
  wire n3604_o;
  wire n3606_o;
  wire n3608_o;
  wire n3610_o;
  wire n3612_o;
  wire [2:0] n3613_o;
  wire [2:0] n3614_o;
  wire n3616_o;
  wire [2:0] n3617_o;
  wire n3619_o;
  wire [1:0] n3620_o;
  wire n3622_o;
  wire n3623_o;
  wire n3624_o;
  wire [1:0] n3625_o;
  wire n3627_o;
  wire n3628_o;
  wire n3629_o;
  wire n3631_o;
  wire n3633_o;
  wire n3634_o;
  wire n3636_o;
  wire n3638_o;
  wire n3639_o;
  wire n3640_o;
  wire n3641_o;
  wire n3643_o;
  wire [1:0] n3644_o;
  wire n3646_o;
  wire n3649_o;
  wire n3650_o;
  wire [1:0] n3652_o;
  wire n3655_o;
  wire n3658_o;
  wire n3661_o;
  wire n3664_o;
  wire n3666_o;
  wire n3668_o;
  wire [1:0] n3672_o;
  wire n3674_o;
  wire n3677_o;
  wire n3679_o;
  wire n3680_o;
  wire n3681_o;
  wire n3682_o;
  wire n3684_o;
  wire n3687_o;
  wire n3689_o;
  wire n3691_o;
  wire n3693_o;
  wire n3694_o;
  wire n3695_o;
  wire n3696_o;
  wire n3697_o;
  wire n3699_o;
  wire n3701_o;
  wire n3703_o;
  wire n3704_o;
  wire n3705_o;
  wire n3706_o;
  wire n3708_o;
  wire n3710_o;
  wire n3713_o;
  wire n3715_o;
  wire n3717_o;
  wire n3719_o;
  wire n3720_o;
  wire n3721_o;
  wire n3722_o;
  wire n3723_o;
  wire [1:0] n3724_o;
  wire [1:0] n3726_o;
  wire n3728_o;
  wire n3730_o;
  wire n3732_o;
  wire [2:0] n3733_o;
  wire n3735_o;
  wire [2:0] n3736_o;
  wire n3738_o;
  wire [1:0] n3739_o;
  wire n3741_o;
  wire n3742_o;
  wire n3743_o;
  wire [1:0] n3744_o;
  wire n3746_o;
  wire n3747_o;
  wire n3749_o;
  wire n3751_o;
  wire [1:0] n3753_o;
  wire n3755_o;
  wire n3758_o;
  wire [1:0] n3760_o;
  wire n3763_o;
  wire n3766_o;
  wire n3769_o;
  wire n3772_o;
  wire n3774_o;
  wire n3776_o;
  wire n3778_o;
  wire n3780_o;
  wire n3781_o;
  wire n3782_o;
  wire n3783_o;
  wire n3785_o;
  wire n3787_o;
  wire n3788_o;
  wire [1:0] n3789_o;
  wire n3791_o;
  wire n3794_o;
  wire n3795_o;
  wire n3796_o;
  wire n3798_o;
  wire n3800_o;
  wire n3802_o;
  wire n3804_o;
  wire n3805_o;
  wire n3806_o;
  wire n3808_o;
  wire n3810_o;
  wire n3811_o;
  wire n3812_o;
  wire n3813_o;
  wire n3815_o;
  wire n3817_o;
  wire n3819_o;
  wire n3821_o;
  wire n3822_o;
  wire n3823_o;
  wire n3825_o;
  wire n3827_o;
  wire n3829_o;
  wire n3831_o;
  wire [1:0] n3832_o;
  wire n3834_o;
  wire [2:0] n3835_o;
  wire n3837_o;
  wire [3:0] n3838_o;
  wire n3840_o;
  wire [1:0] n3841_o;
  wire n3843_o;
  wire n3844_o;
  wire n3845_o;
  wire [1:0] n3846_o;
  wire n3848_o;
  wire n3849_o;
  wire n3851_o;
  wire n3852_o;
  wire n3853_o;
  wire n3854_o;
  wire n3855_o;
  wire n3857_o;
  wire n3858_o;
  wire [1:0] n3860_o;
  wire n3863_o;
  wire n3866_o;
  wire n3869_o;
  wire n3872_o;
  wire n3874_o;
  wire [2:0] n3875_o;
  wire n3877_o;
  wire [2:0] n3878_o;
  wire n3880_o;
  wire [1:0] n3881_o;
  wire n3883_o;
  wire n3884_o;
  wire n3885_o;
  wire [1:0] n3888_o;
  wire n3890_o;
  wire n3893_o;
  wire n3895_o;
  wire n3896_o;
  wire n3899_o;
  wire n3902_o;
  wire n3905_o;
  wire n3908_o;
  wire n3911_o;
  wire n3913_o;
  wire n3914_o;
  wire n3915_o;
  wire n3917_o;
  wire n3919_o;
  wire n3920_o;
  wire n3922_o;
  wire n3923_o;
  wire n3924_o;
  wire n3925_o;
  wire n3926_o;
  wire n3928_o;
  wire n3929_o;
  wire n3930_o;
  wire n3931_o;
  wire n3932_o;
  wire n3934_o;
  wire n3936_o;
  wire n3938_o;
  wire [1:0] n3939_o;
  wire n3941_o;
  wire [2:0] n3942_o;
  wire n3944_o;
  wire [3:0] n3945_o;
  wire n3947_o;
  wire [1:0] n3948_o;
  wire n3950_o;
  wire n3951_o;
  wire n3952_o;
  wire [1:0] n3953_o;
  wire n3955_o;
  wire n3956_o;
  wire n3958_o;
  wire n3959_o;
  wire n3960_o;
  wire n3961_o;
  wire n3962_o;
  wire [1:0] n3965_o;
  wire [1:0] n3966_o;
  wire [1:0] n3967_o;
  wire n3968_o;
  wire [1:0] n3969_o;
  wire n3971_o;
  wire n3972_o;
  wire n3973_o;
  wire n3975_o;
  wire n3976_o;
  wire n3977_o;
  wire n3978_o;
  wire n3979_o;
  wire [1:0] n3981_o;
  wire [1:0] n3983_o;
  wire n3984_o;
  wire n3987_o;
  wire n3990_o;
  wire n3993_o;
  wire n3996_o;
  wire n3998_o;
  wire n3999_o;
  wire n4000_o;
  wire n4002_o;
  wire n4005_o;
  wire n4007_o;
  wire n4009_o;
  wire n4011_o;
  wire n4013_o;
  wire [2:0] n4014_o;
  wire n4016_o;
  wire [2:0] n4017_o;
  wire n4019_o;
  wire [1:0] n4020_o;
  wire n4022_o;
  wire n4023_o;
  wire n4024_o;
  wire [2:0] n4027_o;
  wire n4029_o;
  wire n4032_o;
  wire n4034_o;
  wire n4035_o;
  wire n4038_o;
  wire n4041_o;
  wire n4044_o;
  wire n4047_o;
  wire n4049_o;
  wire n4051_o;
  wire n4053_o;
  wire n4055_o;
  wire n4056_o;
  wire n4057_o;
  wire n4059_o;
  wire n4061_o;
  wire n4062_o;
  wire n4064_o;
  wire n4065_o;
  wire n4066_o;
  wire n4068_o;
  wire n4069_o;
  wire n4070_o;
  wire n4072_o;
  wire n4074_o;
  wire n4076_o;
  wire n4078_o;
  wire n4079_o;
  wire [2:0] n4080_o;
  wire n4082_o;
  wire n4083_o;
  wire n4084_o;
  wire n4085_o;
  wire n4089_o;
  wire n4090_o;
  wire [1:0] n4093_o;
  wire n4095_o;
  wire n4096_o;
  wire n4097_o;
  wire [1:0] n4098_o;
  wire n4100_o;
  wire n4101_o;
  wire [2:0] n4102_o;
  wire n4104_o;
  wire [1:0] n4105_o;
  wire n4107_o;
  wire n4108_o;
  wire n4109_o;
  wire n4110_o;
  wire n4111_o;
  wire n4112_o;
  wire [1:0] n4113_o;
  wire n4115_o;
  wire [2:0] n4116_o;
  wire n4118_o;
  wire n4119_o;
  wire [3:0] n4120_o;
  wire n4122_o;
  wire n4123_o;
  wire n4124_o;
  wire n4125_o;
  wire n4127_o;
  wire n4128_o;
  wire [1:0] n4130_o;
  wire [2:0] n4131_o;
  wire n4133_o;
  wire [2:0] n4134_o;
  wire n4136_o;
  wire n4137_o;
  wire n4139_o;
  wire n4140_o;
  wire n4144_o;
  wire n4146_o;
  wire [2:0] n4147_o;
  wire n4149_o;
  wire n4153_o;
  wire n4154_o;
  wire n4155_o;
  wire n4157_o;
  wire n4158_o;
  wire n4159_o;
  wire n4162_o;
  wire n4163_o;
  wire n4164_o;
  wire n4165_o;
  wire [2:0] n4167_o;
  wire n4169_o;
  wire [2:0] n4170_o;
  wire n4172_o;
  wire n4173_o;
  wire [2:0] n4174_o;
  wire n4176_o;
  wire n4177_o;
  wire n4179_o;
  wire n4180_o;
  wire [6:0] n4183_o;
  wire n4184_o;
  wire n4185_o;
  wire n4186_o;
  wire n4187_o;
  wire [6:0] n4188_o;
  wire n4189_o;
  wire n4191_o;
  wire n4192_o;
  wire [1:0] n4196_o;
  wire n4197_o;
  wire n4198_o;
  wire [1:0] n4201_o;
  wire n4203_o;
  wire n4204_o;
  wire n4205_o;
  wire n4206_o;
  wire n4207_o;
  wire [6:0] n4209_o;
  wire [1:0] n4210_o;
  wire n4212_o;
  wire n4214_o;
  wire n4216_o;
  wire n4217_o;
  wire n4218_o;
  wire n4219_o;
  wire n4222_o;
  wire n4224_o;
  wire n4227_o;
  wire n4230_o;
  wire [1:0] n4231_o;
  wire n4233_o;
  wire n4235_o;
  wire n4237_o;
  wire n4239_o;
  wire [1:0] n4240_o;
  wire n4242_o;
  wire n4244_o;
  wire n4246_o;
  wire n4248_o;
  wire n4250_o;
  wire [6:0] n4251_o;
  wire [1:0] n4252_o;
  wire [1:0] n4253_o;
  wire n4255_o;
  wire n4258_o;
  wire n4260_o;
  wire n4262_o;
  wire n4264_o;
  wire n4265_o;
  wire n4266_o;
  wire n4267_o;
  wire n4268_o;
  wire n4269_o;
  wire n4270_o;
  wire n4271_o;
  wire n4272_o;
  wire [1:0] n4273_o;
  wire n4274_o;
  wire n4275_o;
  wire n4276_o;
  wire n4277_o;
  wire n4278_o;
  wire n4279_o;
  wire n4281_o;
  wire n4283_o;
  wire n4285_o;
  wire n4286_o;
  wire n4288_o;
  wire [6:0] n4289_o;
  wire n4290_o;
  wire [1:0] n4291_o;
  wire n4293_o;
  wire [2:0] n4294_o;
  wire n4296_o;
  wire n4297_o;
  wire [3:0] n4298_o;
  wire n4300_o;
  wire [1:0] n4301_o;
  wire n4303_o;
  wire n4304_o;
  wire n4305_o;
  wire n4307_o;
  wire n4308_o;
  wire n4309_o;
  wire n4310_o;
  wire n4312_o;
  wire n4314_o;
  wire n4315_o;
  wire n4316_o;
  wire n4319_o;
  wire n4320_o;
  wire n4321_o;
  wire n4322_o;
  wire [6:0] n4324_o;
  wire n4326_o;
  wire n4327_o;
  wire [1:0] n4328_o;
  wire n4330_o;
  wire n4331_o;
  wire n4332_o;
  wire n4333_o;
  wire n4336_o;
  wire [1:0] n4338_o;
  wire [6:0] n4340_o;
  wire n4344_o;
  wire n4347_o;
  wire n4348_o;
  wire n4349_o;
  wire n4350_o;
  wire n4351_o;
  wire n4352_o;
  wire n4353_o;
  wire n4354_o;
  wire [1:0] n4355_o;
  wire n4357_o;
  wire [2:0] n4358_o;
  wire n4360_o;
  wire n4361_o;
  wire [3:0] n4362_o;
  wire n4364_o;
  wire [1:0] n4365_o;
  wire n4367_o;
  wire n4368_o;
  wire n4369_o;
  wire n4370_o;
  wire n4371_o;
  wire n4373_o;
  wire n4375_o;
  wire n4376_o;
  wire n4377_o;
  wire n4378_o;
  wire n4379_o;
  wire n4381_o;
  wire n4383_o;
  wire n4384_o;
  wire n4385_o;
  wire n4386_o;
  wire n4389_o;
  wire n4390_o;
  wire n4391_o;
  wire n4392_o;
  wire [6:0] n4394_o;
  wire n4396_o;
  wire n4397_o;
  wire [1:0] n4398_o;
  wire n4400_o;
  wire n4401_o;
  wire n4402_o;
  wire n4403_o;
  wire n4404_o;
  wire n4406_o;
  wire n4407_o;
  wire [6:0] n4410_o;
  wire [1:0] n4412_o;
  wire n4415_o;
  wire n4418_o;
  wire n4419_o;
  wire n4420_o;
  wire [6:0] n4421_o;
  wire [1:0] n4422_o;
  wire n4424_o;
  wire n4425_o;
  wire n4426_o;
  wire n4429_o;
  wire [1:0] n4431_o;
  wire n4432_o;
  wire n4435_o;
  wire n4437_o;
  wire n4439_o;
  wire n4441_o;
  wire n4444_o;
  wire n4447_o;
  wire n4449_o;
  wire n4451_o;
  wire n4453_o;
  wire [6:0] n4454_o;
  wire [1:0] n4456_o;
  wire [1:0] n4457_o;
  wire n4459_o;
  wire n4461_o;
  wire n4462_o;
  wire n4464_o;
  wire n4466_o;
  wire n4468_o;
  wire n4470_o;
  wire n4471_o;
  wire n4472_o;
  wire n4474_o;
  wire n4475_o;
  wire n4477_o;
  wire n4478_o;
  wire [6:0] n4479_o;
  wire n4480_o;
  wire [2:0] n4481_o;
  wire n4483_o;
  wire [2:0] n4486_o;
  wire n4488_o;
  wire n4489_o;
  wire [1:0] n4490_o;
  wire n4492_o;
  wire n4493_o;
  wire [2:0] n4494_o;
  wire n4496_o;
  wire n4497_o;
  wire [3:0] n4498_o;
  wire n4500_o;
  wire n4501_o;
  wire n4503_o;
  wire n4504_o;
  wire [1:0] n4507_o;
  wire n4509_o;
  wire n4510_o;
  wire n4511_o;
  wire n4512_o;
  wire n4513_o;
  wire [6:0] n4515_o;
  wire n4516_o;
  wire [1:0] n4518_o;
  wire [1:0] n4519_o;
  wire n4520_o;
  wire n4523_o;
  wire n4526_o;
  wire n4529_o;
  wire n4532_o;
  wire n4533_o;
  wire n4534_o;
  wire n4535_o;
  wire n4536_o;
  wire n4537_o;
  wire [1:0] n4538_o;
  wire n4539_o;
  wire n4541_o;
  wire n4543_o;
  wire n4545_o;
  wire n4547_o;
  wire n4548_o;
  wire n4549_o;
  wire n4550_o;
  wire n4551_o;
  wire [6:0] n4552_o;
  wire [1:0] n4553_o;
  wire n4554_o;
  wire n4556_o;
  wire n4558_o;
  wire n4560_o;
  wire n4562_o;
  wire n4563_o;
  wire n4564_o;
  wire n4565_o;
  wire n4566_o;
  wire n4568_o;
  wire n4570_o;
  wire [6:0] n4571_o;
  wire [2:0] n4572_o;
  wire n4574_o;
  wire n4584_o;
  wire n4587_o;
  wire n4590_o;
  wire n4591_o;
  wire n4592_o;
  wire n4593_o;
  wire n4594_o;
  wire n4595_o;
  wire n4596_o;
  wire n4597_o;
  wire n4598_o;
  wire n4599_o;
  wire n4600_o;
  wire n4601_o;
  wire [6:0] n4603_o;
  wire [2:0] n4604_o;
  wire n4606_o;
  wire [2:0] n4607_o;
  wire n4609_o;
  wire [1:0] n4610_o;
  wire n4612_o;
  wire n4613_o;
  wire n4614_o;
  wire [1:0] n4619_o;
  wire n4621_o;
  wire n4624_o;
  wire n4626_o;
  wire n4627_o;
  wire n4630_o;
  wire n4633_o;
  wire n4636_o;
  wire n4639_o;
  wire n4642_o;
  wire n4644_o;
  wire n4645_o;
  wire n4646_o;
  wire n4648_o;
  wire n4650_o;
  wire n4652_o;
  wire n4654_o;
  wire [1:0] n4656_o;
  wire n4658_o;
  wire n4659_o;
  wire n4661_o;
  wire n4662_o;
  wire n4664_o;
  wire n4666_o;
  wire n4668_o;
  wire n4670_o;
  wire n4672_o;
  wire n4673_o;
  wire n4674_o;
  wire n4675_o;
  wire n4676_o;
  wire n4677_o;
  wire n4678_o;
  wire n4679_o;
  wire n4680_o;
  wire n4682_o;
  wire n4683_o;
  wire n4684_o;
  wire n4685_o;
  wire n4686_o;
  wire n4688_o;
  wire n4690_o;
  wire n4691_o;
  wire n4692_o;
  wire [1:0] n4694_o;
  wire [1:0] n4695_o;
  wire n4697_o;
  wire n4698_o;
  wire n4700_o;
  wire n4702_o;
  wire n4704_o;
  wire n4705_o;
  wire n4706_o;
  wire n4707_o;
  wire [2:0] n4708_o;
  wire n4709_o;
  wire n4710_o;
  wire n4711_o;
  wire n4712_o;
  wire n4713_o;
  wire n4714_o;
  wire n4715_o;
  wire [2:0] n4716_o;
  wire [2:0] n4717_o;
  wire n4718_o;
  wire n4720_o;
  wire n4722_o;
  wire n4724_o;
  wire n4726_o;
  wire n4727_o;
  wire [6:0] n4728_o;
  wire [1:0] n4729_o;
  wire [1:0] n4730_o;
  wire n4732_o;
  wire n4733_o;
  wire n4735_o;
  wire n4737_o;
  wire n4738_o;
  wire n4740_o;
  wire n4742_o;
  wire n4744_o;
  wire n4745_o;
  wire n4746_o;
  wire n4748_o;
  wire n4750_o;
  wire n4751_o;
  wire n4752_o;
  wire n4754_o;
  wire n4755_o;
  wire n4756_o;
  wire n4757_o;
  wire n4758_o;
  wire n4759_o;
  wire n4760_o;
  wire n4761_o;
  wire n4762_o;
  wire n4763_o;
  wire n4764_o;
  wire n4765_o;
  wire n4766_o;
  wire [2:0] n4767_o;
  wire [2:0] n4768_o;
  wire n4770_o;
  wire n4771_o;
  wire n4772_o;
  wire n4773_o;
  wire n4775_o;
  wire n4777_o;
  wire n4779_o;
  wire n4781_o;
  wire n4783_o;
  wire [6:0] n4784_o;
  wire [1:0] n4785_o;
  wire [1:0] n4786_o;
  wire n4788_o;
  wire n4789_o;
  wire n4790_o;
  wire n4792_o;
  wire n4793_o;
  wire n4795_o;
  wire n4797_o;
  wire n4799_o;
  wire n4801_o;
  wire n4802_o;
  wire n4803_o;
  wire n4805_o;
  wire n4806_o;
  wire n4807_o;
  wire n4808_o;
  wire n4809_o;
  wire n4810_o;
  wire n4811_o;
  wire n4812_o;
  wire n4813_o;
  wire n4814_o;
  wire n4815_o;
  wire n4816_o;
  wire n4817_o;
  wire n4818_o;
  wire n4819_o;
  wire n4820_o;
  wire n4821_o;
  wire n4822_o;
  wire n4823_o;
  wire n4824_o;
  wire n4825_o;
  wire n4826_o;
  wire n4827_o;
  wire n4828_o;
  wire n4829_o;
  wire n4830_o;
  wire n4831_o;
  wire n4832_o;
  wire n4833_o;
  wire n4834_o;
  wire n4835_o;
  wire n4836_o;
  wire n4837_o;
  wire n4838_o;
  wire n4839_o;
  wire n4840_o;
  wire n4841_o;
  wire n4842_o;
  wire n4844_o;
  wire n4846_o;
  wire n4848_o;
  wire n4850_o;
  wire n4852_o;
  wire n4854_o;
  wire n4856_o;
  wire n4857_o;
  wire n4859_o;
  wire [6:0] n4860_o;
  wire n4862_o;
  wire n4864_o;
  wire n4865_o;
  wire [4:0] n4866_o;
  wire n4868_o;
  wire [1:0] n4869_o;
  wire n4871_o;
  wire n4872_o;
  wire [1:0] n4873_o;
  wire n4875_o;
  wire [2:0] n4876_o;
  wire n4878_o;
  wire [2:0] n4879_o;
  wire n4881_o;
  wire [1:0] n4882_o;
  wire n4884_o;
  wire n4885_o;
  wire n4886_o;
  wire n4887_o;
  wire [1:0] n4888_o;
  wire n4890_o;
  wire [2:0] n4891_o;
  wire n4893_o;
  wire n4894_o;
  wire [3:0] n4895_o;
  wire n4897_o;
  wire [1:0] n4898_o;
  wire n4900_o;
  wire n4901_o;
  wire n4902_o;
  wire n4903_o;
  wire n4904_o;
  wire n4907_o;
  wire n4909_o;
  wire n4912_o;
  wire [1:0] n4914_o;
  wire n4916_o;
  wire [1:0] n4917_o;
  wire n4919_o;
  wire n4922_o;
  wire [1:0] n4924_o;
  wire n4927_o;
  wire n4930_o;
  wire n4932_o;
  wire n4933_o;
  wire n4935_o;
  wire n4937_o;
  wire n4939_o;
  wire n4941_o;
  wire n4944_o;
  wire n4947_o;
  wire n4950_o;
  wire n4952_o;
  wire n4954_o;
  wire [1:0] n4955_o;
  wire n4957_o;
  wire n4959_o;
  wire n4961_o;
  wire n4963_o;
  wire n4965_o;
  wire n4967_o;
  wire n4969_o;
  wire n4971_o;
  wire n4973_o;
  wire n4975_o;
  wire n4976_o;
  wire n4977_o;
  wire [1:0] n4978_o;
  wire n4980_o;
  wire n4981_o;
  wire [2:0] n4982_o;
  wire n4984_o;
  wire n4985_o;
  wire [3:0] n4986_o;
  wire n4988_o;
  wire n4989_o;
  wire n4990_o;
  wire [6:0] n4992_o;
  wire n4994_o;
  wire n4995_o;
  wire n4996_o;
  wire n4997_o;
  wire n4998_o;
  wire [1:0] n5001_o;
  wire n5003_o;
  wire n5004_o;
  wire n5005_o;
  wire n5006_o;
  wire n5007_o;
  wire [6:0] n5009_o;
  wire n5011_o;
  wire n5012_o;
  wire n5013_o;
  wire n5014_o;
  wire n5016_o;
  wire n5018_o;
  wire n5021_o;
  wire n5023_o;
  wire n5024_o;
  wire n5025_o;
  wire n5026_o;
  wire n5028_o;
  wire n5030_o;
  wire [1:0] n5032_o;
  wire n5033_o;
  wire n5034_o;
  wire n5035_o;
  wire [1:0] n5037_o;
  wire [1:0] n5038_o;
  wire n5039_o;
  wire n5041_o;
  wire n5044_o;
  wire n5047_o;
  wire n5050_o;
  wire n5053_o;
  wire [1:0] n5054_o;
  wire n5055_o;
  wire n5056_o;
  wire n5057_o;
  wire n5058_o;
  wire [1:0] n5059_o;
  wire [6:0] n5060_o;
  wire [6:0] n5061_o;
  wire n5063_o;
  wire n5065_o;
  wire n5066_o;
  wire n5068_o;
  wire n5069_o;
  wire n5071_o;
  wire n5072_o;
  wire n5074_o;
  wire n5075_o;
  wire n5077_o;
  wire n5078_o;
  wire n5080_o;
  wire n5081_o;
  wire n5083_o;
  wire n5084_o;
  wire n5086_o;
  wire n5087_o;
  wire n5089_o;
  wire n5090_o;
  wire n5092_o;
  wire n5093_o;
  wire n5095_o;
  wire n5096_o;
  wire n5098_o;
  wire n5099_o;
  wire n5101_o;
  wire n5102_o;
  wire n5104_o;
  wire n5105_o;
  wire n5107_o;
  wire n5108_o;
  wire n5116_o;
  wire n5119_o;
  wire n5122_o;
  wire n5123_o;
  wire n5124_o;
  wire n5125_o;
  wire n5126_o;
  wire n5127_o;
  wire n5128_o;
  wire n5129_o;
  wire n5130_o;
  wire [6:0] n5132_o;
  wire n5134_o;
  wire n5136_o;
  wire n5137_o;
  wire n5139_o;
  wire n5140_o;
  wire n5142_o;
  wire n5143_o;
  wire n5145_o;
  wire n5146_o;
  wire n5148_o;
  wire n5149_o;
  wire n5151_o;
  wire n5152_o;
  wire n5154_o;
  wire n5155_o;
  wire [1:0] n5162_o;
  wire n5164_o;
  wire n5167_o;
  wire n5170_o;
  wire n5171_o;
  wire n5172_o;
  wire n5173_o;
  wire n5174_o;
  wire [6:0] n5176_o;
  wire n5178_o;
  wire n5180_o;
  wire n5181_o;
  wire n5183_o;
  wire n5184_o;
  wire n5186_o;
  wire n5187_o;
  wire n5189_o;
  wire n5190_o;
  wire n5192_o;
  wire n5193_o;
  wire n5195_o;
  wire n5196_o;
  wire n5198_o;
  wire n5199_o;
  wire [1:0] n5202_o;
  wire n5205_o;
  wire n5208_o;
  wire n5211_o;
  wire n5214_o;
  wire n5215_o;
  wire n5216_o;
  wire n5217_o;
  wire n5218_o;
  wire n5220_o;
  wire n5222_o;
  wire n5223_o;
  wire n5225_o;
  wire n5226_o;
  wire n5228_o;
  wire n5229_o;
  wire n5231_o;
  wire n5232_o;
  wire n5234_o;
  wire n5235_o;
  wire n5237_o;
  wire n5238_o;
  wire n5240_o;
  wire n5241_o;
  wire [1:0] n5245_o;
  wire n5248_o;
  wire n5251_o;
  wire n5252_o;
  wire n5253_o;
  wire n5254_o;
  wire n5255_o;
  wire n5257_o;
  wire n5259_o;
  wire n5261_o;
  wire n5262_o;
  wire n5264_o;
  wire n5265_o;
  wire n5267_o;
  wire n5268_o;
  wire n5270_o;
  wire n5271_o;
  wire n5273_o;
  wire n5274_o;
  wire n5276_o;
  wire n5277_o;
  wire n5279_o;
  wire n5280_o;
  wire n5281_o;
  wire [5:0] n5285_o;
  wire n5286_o;
  wire n5287_o;
  wire [5:0] n5288_o;
  wire n5291_o;
  wire n5294_o;
  wire n5295_o;
  wire n5296_o;
  wire n5297_o;
  wire n5298_o;
  wire n5300_o;
  wire n5302_o;
  wire n5303_o;
  wire n5305_o;
  wire n5308_o;
  wire n5310_o;
  wire n5311_o;
  wire n5312_o;
  wire n5315_o;
  wire n5318_o;
  wire n5320_o;
  wire n5322_o;
  wire n5323_o;
  wire n5324_o;
  wire n5326_o;
  wire n5329_o;
  wire n5330_o;
  wire n5331_o;
  wire n5332_o;
  wire [1:0] n5334_o;
  wire n5336_o;
  wire [1:0] n5337_o;
  wire n5338_o;
  wire n5339_o;
  wire n5340_o;
  wire n5341_o;
  wire [1:0] n5342_o;
  wire [1:0] n5343_o;
  wire [6:0] n5345_o;
  wire n5346_o;
  wire n5347_o;
  wire n5350_o;
  wire n5353_o;
  wire n5354_o;
  wire n5355_o;
  wire n5356_o;
  wire n5357_o;
  wire n5359_o;
  wire n5360_o;
  wire n5362_o;
  wire n5364_o;
  wire n5365_o;
  wire [1:0] n5370_o;
  wire n5372_o;
  wire n5374_o;
  wire [1:0] n5375_o;
  wire n5376_o;
  wire n5377_o;
  wire n5378_o;
  wire n5379_o;
  wire [1:0] n5380_o;
  wire [1:0] n5381_o;
  wire [6:0] n5383_o;
  wire n5385_o;
  wire [1:0] n5390_o;
  wire n5392_o;
  wire [1:0] n5393_o;
  wire n5394_o;
  wire n5395_o;
  wire n5396_o;
  wire n5397_o;
  wire [1:0] n5398_o;
  wire [1:0] n5399_o;
  wire [6:0] n5401_o;
  wire n5403_o;
  wire [1:0] n5405_o;
  wire n5406_o;
  wire n5408_o;
  wire n5409_o;
  wire n5412_o;
  wire n5415_o;
  wire n5417_o;
  wire n5419_o;
  wire n5420_o;
  wire [11:0] n5421_o;
  wire n5423_o;
  wire n5425_o;
  wire n5427_o;
  wire n5428_o;
  wire n5429_o;
  wire n5430_o;
  wire [1:0] n5431_o;
  wire [1:0] n5432_o;
  wire n5433_o;
  wire n5434_o;
  wire n5438_o;
  wire n5440_o;
  wire n5442_o;
  wire [6:0] n5444_o;
  wire [1:0] n5446_o;
  wire n5447_o;
  wire n5450_o;
  wire n5453_o;
  wire [1:0] n5454_o;
  wire [1:0] n5455_o;
  wire [1:0] n5457_o;
  wire [6:0] n5458_o;
  wire [1:0] n5459_o;
  wire n5460_o;
  wire n5463_o;
  wire n5465_o;
  wire n5467_o;
  wire [1:0] n5468_o;
  wire [1:0] n5470_o;
  wire [6:0] n5471_o;
  wire n5473_o;
  wire n5475_o;
  wire n5476_o;
  wire [12:0] n5477_o;
  reg n5478_o;
  reg [1:0] n5483_o;
  reg [1:0] n5484_o;
  reg n5485_o;
  reg n5486_o;
  reg n5487_o;
  reg n5489_o;
  reg n5491_o;
  reg [5:0] n5492_o;
  reg n5493_o;
  reg n5496_o;
  reg n5498_o;
  reg n5501_o;
  reg n5503_o;
  reg n5507_o;
  reg n5509_o;
  wire n5510_o;
  reg n5511_o;
  wire n5512_o;
  reg n5513_o;
  wire n5514_o;
  reg n5515_o;
  wire n5516_o;
  reg n5517_o;
  wire n5518_o;
  wire n5519_o;
  wire n5520_o;
  reg n5521_o;
  wire n5522_o;
  wire n5523_o;
  wire n5524_o;
  reg n5525_o;
  wire n5526_o;
  reg n5527_o;
  wire n5528_o;
  reg n5529_o;
  wire [1:0] n5530_o;
  reg [1:0] n5531_o;
  wire [1:0] n5532_o;
  reg [1:0] n5533_o;
  wire n5534_o;
  wire n5535_o;
  wire n5536_o;
  wire n5537_o;
  reg n5538_o;
  wire n5539_o;
  wire n5540_o;
  wire n5541_o;
  wire n5542_o;
  reg n5543_o;
  wire n5544_o;
  reg n5545_o;
  reg n5547_o;
  reg n5549_o;
  reg [1:0] n5551_o;
  reg n5553_o;
  reg [6:0] n5554_o;
  wire n5555_o;
  wire [1:0] n5556_o;
  wire [1:0] n5557_o;
  wire n5558_o;
  wire n5559_o;
  wire n5560_o;
  wire n5562_o;
  wire n5564_o;
  wire n5566_o;
  wire n5568_o;
  wire [5:0] n5569_o;
  wire n5570_o;
  wire n5571_o;
  wire n5573_o;
  wire n5575_o;
  wire n5577_o;
  wire n5578_o;
  wire n5580_o;
  wire n5582_o;
  wire [1:0] n5583_o;
  wire [3:0] n5584_o;
  wire [1:0] n5585_o;
  wire n5586_o;
  wire n5587_o;
  wire n5588_o;
  wire n5589_o;
  wire n5590_o;
  wire n5591_o;
  wire n5592_o;
  wire n5593_o;
  wire n5594_o;
  wire n5595_o;
  wire n5596_o;
  wire n5597_o;
  wire n5598_o;
  wire n5599_o;
  wire n5600_o;
  wire n5601_o;
  wire n5602_o;
  wire n5603_o;
  wire n5604_o;
  wire [3:0] n5605_o;
  wire [3:0] n5606_o;
  wire n5607_o;
  wire [1:0] n5608_o;
  wire n5609_o;
  wire n5610_o;
  wire [2:0] n5611_o;
  wire n5613_o;
  wire n5615_o;
  wire [2:0] n5617_o;
  wire [6:0] n5618_o;
  wire n5620_o;
  wire [6:0] n5621_o;
  reg n5622_o;
  reg [1:0] n5623_o;
  reg [1:0] n5624_o;
  reg n5625_o;
  reg n5626_o;
  reg n5628_o;
  reg n5629_o;
  reg n5631_o;
  reg n5633_o;
  reg n5635_o;
  reg n5637_o;
  reg n5639_o;
  reg n5641_o;
  reg n5643_o;
  reg n5645_o;
  reg [5:0] n5646_o;
  reg n5648_o;
  reg n5649_o;
  reg n5651_o;
  reg n5653_o;
  reg n5655_o;
  reg n5657_o;
  reg n5659_o;
  reg n5661_o;
  reg n5663_o;
  wire n5664_o;
  reg n5665_o;
  wire n5666_o;
  reg n5667_o;
  wire n5668_o;
  reg n5669_o;
  wire n5670_o;
  reg n5671_o;
  wire n5672_o;
  reg n5673_o;
  wire n5674_o;
  reg n5675_o;
  wire n5676_o;
  reg n5677_o;
  wire n5678_o;
  reg n5679_o;
  wire n5680_o;
  wire n5681_o;
  wire n5682_o;
  reg n5683_o;
  wire n5684_o;
  wire n5685_o;
  wire n5686_o;
  reg n5687_o;
  wire n5688_o;
  reg n5689_o;
  wire n5690_o;
  reg n5691_o;
  wire n5692_o;
  wire n5693_o;
  reg n5694_o;
  wire n5695_o;
  wire n5696_o;
  reg n5697_o;
  wire n5698_o;
  reg n5699_o;
  wire n5700_o;
  reg n5701_o;
  wire n5702_o;
  reg n5703_o;
  wire n5704_o;
  reg n5705_o;
  wire [3:0] n5706_o;
  reg [3:0] n5707_o;
  reg [1:0] n5708_o;
  reg [1:0] n5709_o;
  wire n5710_o;
  reg n5711_o;
  wire n5712_o;
  reg n5713_o;
  wire n5714_o;
  reg n5715_o;
  reg n5716_o;
  wire n5717_o;
  reg n5718_o;
  reg n5720_o;
  wire n5721_o;
  reg n5723_o;
  wire n5724_o;
  reg n5726_o;
  reg n5728_o;
  reg n5730_o;
  reg n5732_o;
  reg n5734_o;
  reg n5736_o;
  reg n5738_o;
  reg n5740_o;
  reg n5742_o;
  wire [1:0] n5743_o;
  reg [1:0] n5745_o;
  wire n5746_o;
  reg n5748_o;
  reg n5750_o;
  reg [6:0] n5751_o;
  wire n5752_o;
  wire [1:0] n5753_o;
  wire [1:0] n5754_o;
  wire n5755_o;
  wire n5756_o;
  wire n5758_o;
  wire n5759_o;
  wire n5761_o;
  wire n5763_o;
  wire n5764_o;
  wire n5765_o;
  wire n5766_o;
  wire n5768_o;
  wire n5770_o;
  wire n5772_o;
  wire n5773_o;
  wire [5:0] n5774_o;
  wire n5776_o;
  wire n5777_o;
  wire n5778_o;
  wire n5780_o;
  wire n5782_o;
  wire n5784_o;
  wire n5785_o;
  wire n5787_o;
  wire n5788_o;
  wire [3:0] n5789_o;
  wire [9:0] n5790_o;
  wire [4:0] n5791_o;
  wire [1:0] n5792_o;
  wire n5793_o;
  wire n5794_o;
  wire n5795_o;
  wire n5796_o;
  wire n5797_o;
  wire n5798_o;
  wire n5799_o;
  wire n5800_o;
  wire n5801_o;
  wire n5802_o;
  wire n5803_o;
  wire n5804_o;
  wire n5805_o;
  wire n5806_o;
  wire n5807_o;
  wire n5808_o;
  wire n5809_o;
  wire n5810_o;
  wire [2:0] n5811_o;
  wire n5812_o;
  wire [2:0] n5813_o;
  wire [2:0] n5814_o;
  wire n5815_o;
  wire n5816_o;
  wire [4:0] n5817_o;
  wire [4:0] n5818_o;
  wire [4:0] n5819_o;
  wire n5820_o;
  wire n5821_o;
  wire [3:0] n5822_o;
  wire [3:0] n5823_o;
  wire [3:0] n5824_o;
  wire n5825_o;
  wire [4:0] n5826_o;
  wire [4:0] n5827_o;
  wire n5828_o;
  wire n5829_o;
  wire n5830_o;
  wire n5831_o;
  wire n5832_o;
  wire [1:0] n5833_o;
  wire [1:0] n5834_o;
  wire [1:0] n5835_o;
  wire [1:0] n5836_o;
  wire [2:0] n5837_o;
  wire n5838_o;
  wire [1:0] n5840_o;
  wire [1:0] n5842_o;
  wire n5843_o;
  wire n5845_o;
  wire n5847_o;
  wire n5849_o;
  wire n5851_o;
  wire n5853_o;
  wire n5855_o;
  wire [1:0] n5856_o;
  wire [1:0] n5858_o;
  wire n5859_o;
  wire n5860_o;
  wire n5861_o;
  wire [6:0] n5862_o;
  wire n5864_o;
  wire [1:0] n5865_o;
  wire n5867_o;
  wire [2:0] n5868_o;
  wire n5870_o;
  wire n5874_o;
  wire n5875_o;
  wire n5876_o;
  wire [6:0] n5878_o;
  wire [2:0] n5879_o;
  wire n5881_o;
  wire [1:0] n5882_o;
  wire n5884_o;
  wire [2:0] n5885_o;
  wire n5887_o;
  wire n5888_o;
  wire n5889_o;
  wire n5890_o;
  wire [1:0] n5891_o;
  wire n5893_o;
  wire n5894_o;
  wire n5896_o;
  wire n5897_o;
  wire [6:0] n5899_o;
  wire [1:0] n5901_o;
  wire [1:0] n5902_o;
  wire n5903_o;
  wire n5904_o;
  wire n5905_o;
  wire n5906_o;
  wire n5909_o;
  wire n5912_o;
  wire [1:0] n5913_o;
  wire n5916_o;
  wire n5918_o;
  wire n5920_o;
  wire n5921_o;
  wire n5922_o;
  wire [2:0] n5923_o;
  wire n5925_o;
  wire [1:0] n5926_o;
  wire n5928_o;
  wire n5929_o;
  wire n5931_o;
  wire n5933_o;
  wire n5934_o;
  wire n5935_o;
  wire n5936_o;
  wire n5938_o;
  wire [1:0] n5939_o;
  wire n5941_o;
  wire n5944_o;
  wire n5945_o;
  wire [1:0] n5947_o;
  wire n5950_o;
  wire n5953_o;
  wire n5956_o;
  wire n5959_o;
  wire n5961_o;
  wire n5963_o;
  wire n5964_o;
  wire [1:0] n5965_o;
  wire n5966_o;
  wire n5968_o;
  wire n5969_o;
  wire n5971_o;
  wire n5972_o;
  wire n5974_o;
  wire n5975_o;
  wire n5977_o;
  wire n5979_o;
  wire n5980_o;
  wire n5981_o;
  wire [1:0] n5982_o;
  wire [1:0] n5983_o;
  wire n5985_o;
  wire n5987_o;
  wire n5989_o;
  wire n5991_o;
  wire n5993_o;
  wire n5995_o;
  wire n5997_o;
  wire n5998_o;
  wire n6000_o;
  wire n6002_o;
  wire [6:0] n6003_o;
  wire [4:0] n6004_o;
  wire n6006_o;
  wire [2:0] n6007_o;
  wire n6009_o;
  wire [1:0] n6010_o;
  wire n6012_o;
  wire n6013_o;
  wire n6014_o;
  wire [2:0] n6015_o;
  wire n6017_o;
  wire n6019_o;
  wire n6020_o;
  wire n6021_o;
  wire n6023_o;
  wire n6024_o;
  wire [1:0] n6028_o;
  wire n6030_o;
  wire n6033_o;
  wire n6036_o;
  wire n6039_o;
  wire n6042_o;
  wire n6045_o;
  wire n6047_o;
  wire n6049_o;
  wire [1:0] n6050_o;
  wire [1:0] n6052_o;
  wire n6054_o;
  wire n6056_o;
  wire n6057_o;
  wire [1:0] n6058_o;
  wire [1:0] n6059_o;
  wire n6061_o;
  wire n6062_o;
  wire n6063_o;
  wire n6065_o;
  wire n6066_o;
  wire n6067_o;
  wire n6068_o;
  wire n6069_o;
  wire n6071_o;
  wire n6072_o;
  wire n6073_o;
  wire n6074_o;
  wire [1:0] n6076_o;
  wire n6078_o;
  wire n6080_o;
  wire n6081_o;
  wire [6:0] n6082_o;
  wire n6084_o;
  wire n6086_o;
  wire [3:0] n6087_o;
  wire n6089_o;
  wire [7:0] n6091_o;
  wire n6093_o;
  wire [7:0] n6095_o;
  wire n6097_o;
  wire [1:0] n6099_o;
  wire n6102_o;
  wire [6:0] n6105_o;
  wire [1:0] n6106_o;
  wire n6108_o;
  wire n6109_o;
  wire [6:0] n6111_o;
  wire [7:0] n6112_o;
  wire n6114_o;
  wire [7:0] n6116_o;
  wire n6118_o;
  wire [1:0] n6120_o;
  wire [1:0] n6121_o;
  wire n6122_o;
  wire [1:0] n6123_o;
  wire n6125_o;
  wire n6127_o;
  wire n6128_o;
  wire n6129_o;
  wire n6130_o;
  wire n6131_o;
  wire n6132_o;
  wire [6:0] n6134_o;
  wire [1:0] n6135_o;
  wire n6136_o;
  wire n6138_o;
  wire n6139_o;
  wire n6140_o;
  wire n6141_o;
  wire n6142_o;
  wire n6143_o;
  wire [6:0] n6144_o;
  wire n6146_o;
  wire n6147_o;
  wire n6148_o;
  wire [1:0] n6153_o;
  wire n6156_o;
  wire n6159_o;
  wire n6162_o;
  wire [1:0] n6163_o;
  wire [1:0] n6165_o;
  wire n6167_o;
  wire n6169_o;
  wire [1:0] n6170_o;
  wire n6172_o;
  wire [2:0] n6173_o;
  wire n6175_o;
  wire n6177_o;
  wire [3:0] n6178_o;
  wire n6180_o;
  wire [1:0] n6181_o;
  wire n6183_o;
  wire n6184_o;
  wire n6185_o;
  wire [1:0] n6186_o;
  wire n6188_o;
  wire n6191_o;
  wire n6193_o;
  wire n6194_o;
  wire [1:0] n6195_o;
  wire n6197_o;
  wire n6198_o;
  wire n6199_o;
  wire [1:0] n6201_o;
  wire [6:0] n6203_o;
  wire n6204_o;
  wire n6205_o;
  wire n6206_o;
  wire n6209_o;
  wire [1:0] n6210_o;
  wire n6212_o;
  wire n6213_o;
  wire n6214_o;
  wire n6217_o;
  wire [1:0] n6219_o;
  wire n6220_o;
  wire n6222_o;
  wire n6225_o;
  wire n6227_o;
  wire n6230_o;
  wire n6233_o;
  wire n6236_o;
  wire n6238_o;
  wire n6239_o;
  wire n6240_o;
  wire [1:0] n6241_o;
  wire n6243_o;
  wire n6244_o;
  wire [1:0] n6245_o;
  wire n6247_o;
  wire [1:0] n6251_o;
  wire n6253_o;
  wire [1:0] n6254_o;
  wire n6256_o;
  wire n6257_o;
  wire [1:0] n6260_o;
  wire n6262_o;
  wire [1:0] n6267_o;
  wire n6269_o;
  wire n6271_o;
  wire n6272_o;
  wire n6273_o;
  wire [1:0] n6274_o;
  wire n6276_o;
  wire [1:0] n6279_o;
  wire n6283_o;
  wire n6284_o;
  wire n6285_o;
  wire n6286_o;
  wire [6:0] n6288_o;
  wire n6290_o;
  wire [6:0] n6292_o;
  wire [1:0] n6293_o;
  wire n6296_o;
  wire n6299_o;
  wire n6300_o;
  wire n6302_o;
  wire n6304_o;
  wire n6306_o;
  wire [6:0] n6307_o;
  wire [1:0] n6308_o;
  wire n6309_o;
  wire n6311_o;
  wire n6314_o;
  wire n6316_o;
  wire n6317_o;
  wire n6320_o;
  wire n6323_o;
  wire n6325_o;
  wire n6326_o;
  wire n6327_o;
  wire n6329_o;
  wire [1:0] n6330_o;
  wire n6332_o;
  wire n6334_o;
  wire [1:0] n6336_o;
  wire [6:0] n6337_o;
  wire [1:0] n6338_o;
  wire [1:0] n6339_o;
  wire n6341_o;
  wire n6343_o;
  wire n6345_o;
  wire n6346_o;
  wire n6348_o;
  wire n6350_o;
  wire n6353_o;
  wire n6354_o;
  wire n6355_o;
  wire n6356_o;
  wire n6357_o;
  wire n6358_o;
  wire n6359_o;
  wire n6360_o;
  wire n6361_o;
  wire n6363_o;
  wire n6365_o;
  wire n6367_o;
  wire n6369_o;
  wire [1:0] n6371_o;
  wire [6:0] n6372_o;
  wire [1:0] n6373_o;
  wire n6375_o;
  wire n6376_o;
  wire n6377_o;
  wire [2:0] n6378_o;
  wire n6380_o;
  wire n6381_o;
  wire [3:0] n6382_o;
  wire n6384_o;
  wire [1:0] n6385_o;
  wire n6387_o;
  wire n6388_o;
  wire n6389_o;
  wire n6390_o;
  wire [1:0] n6391_o;
  wire n6393_o;
  wire n6394_o;
  wire [2:0] n6395_o;
  wire n6397_o;
  wire [1:0] n6398_o;
  wire n6400_o;
  wire n6401_o;
  wire n6402_o;
  wire n6403_o;
  wire n6404_o;
  wire n6408_o;
  wire n6411_o;
  wire n6414_o;
  wire n6416_o;
  wire [1:0] n6417_o;
  wire [1:0] n6418_o;
  wire n6420_o;
  wire n6422_o;
  wire n6424_o;
  wire n6425_o;
  wire n6426_o;
  wire n6427_o;
  wire n6429_o;
  wire n6431_o;
  wire n6432_o;
  wire n6433_o;
  wire n6434_o;
  wire n6435_o;
  wire n6437_o;
  wire n6438_o;
  wire n6439_o;
  wire n6441_o;
  wire n6443_o;
  wire n6445_o;
  wire n6447_o;
  wire n6449_o;
  wire [1:0] n6451_o;
  wire [6:0] n6452_o;
  wire [1:0] n6453_o;
  wire [1:0] n6454_o;
  wire n6455_o;
  wire n6457_o;
  wire n6459_o;
  wire n6460_o;
  wire n6461_o;
  wire n6462_o;
  wire n6463_o;
  wire n6464_o;
  wire n6466_o;
  wire n6468_o;
  wire n6470_o;
  wire n6471_o;
  wire n6472_o;
  wire n6473_o;
  wire n6474_o;
  wire n6475_o;
  wire n6476_o;
  wire n6477_o;
  wire n6478_o;
  wire n6480_o;
  wire n6482_o;
  wire n6484_o;
  wire n6486_o;
  wire n6487_o;
  wire [1:0] n6489_o;
  wire [6:0] n6490_o;
  wire n6492_o;
  wire [5:0] n6493_o;
  wire n6495_o;
  wire n6496_o;
  wire n6497_o;
  wire [1:0] n6498_o;
  wire n6500_o;
  wire n6501_o;
  wire [3:0] n6502_o;
  wire n6504_o;
  wire [1:0] n6505_o;
  wire n6507_o;
  wire n6508_o;
  wire n6509_o;
  wire n6510_o;
  wire [2:0] n6511_o;
  wire n6513_o;
  wire [1:0] n6514_o;
  wire n6516_o;
  wire n6517_o;
  wire n6518_o;
  wire n6519_o;
  wire n6520_o;
  wire n6522_o;
  wire n6523_o;
  wire n6525_o;
  wire n6526_o;
  wire [1:0] n6527_o;
  wire n6529_o;
  wire n6530_o;
  wire n6531_o;
  wire [1:0] n6533_o;
  wire n6535_o;
  wire n6538_o;
  wire n6542_o;
  wire n6545_o;
  wire n6546_o;
  wire [1:0] n6547_o;
  wire n6549_o;
  wire n6550_o;
  wire n6553_o;
  wire n6556_o;
  wire n6557_o;
  wire n6559_o;
  wire n6562_o;
  wire n6564_o;
  wire n6566_o;
  wire n6568_o;
  wire n6570_o;
  wire n6571_o;
  wire n6572_o;
  wire n6574_o;
  wire n6575_o;
  wire n6577_o;
  wire n6579_o;
  wire n6581_o;
  wire n6583_o;
  wire n6586_o;
  wire n6589_o;
  wire n6592_o;
  wire n6594_o;
  wire n6596_o;
  wire n6598_o;
  wire n6600_o;
  wire n6602_o;
  wire n6604_o;
  wire n6606_o;
  wire n6608_o;
  wire n6609_o;
  wire n6611_o;
  wire [1:0] n6612_o;
  wire n6614_o;
  wire [3:0] n6615_o;
  wire n6617_o;
  wire [1:0] n6618_o;
  wire n6620_o;
  wire n6621_o;
  wire n6622_o;
  wire n6623_o;
  wire [1:0] n6626_o;
  wire n6628_o;
  wire n6630_o;
  wire n6633_o;
  wire n6635_o;
  wire n6638_o;
  wire n6641_o;
  wire n6644_o;
  wire n6646_o;
  wire n6648_o;
  wire n6650_o;
  wire n6652_o;
  wire n6654_o;
  wire n6657_o;
  wire n6660_o;
  wire n6663_o;
  wire n6664_o;
  wire n6665_o;
  wire n6667_o;
  wire n6669_o;
  wire n6670_o;
  wire [2:0] n6671_o;
  wire n6673_o;
  wire [2:0] n6675_o;
  wire n6677_o;
  wire n6679_o;
  wire [1:0] n6683_o;
  wire n6684_o;
  wire n6685_o;
  wire n6686_o;
  wire n6687_o;
  wire n6688_o;
  wire n6689_o;
  wire [6:0] n6691_o;
  wire [2:0] n6694_o;
  wire n6696_o;
  wire [1:0] n6697_o;
  wire n6699_o;
  wire n6700_o;
  wire n6704_o;
  wire n6707_o;
  wire n6710_o;
  wire n6713_o;
  wire n6715_o;
  wire n6716_o;
  wire n6718_o;
  wire n6720_o;
  wire n6722_o;
  wire n6724_o;
  wire n6725_o;
  wire n6726_o;
  wire n6727_o;
  wire n6728_o;
  wire n6729_o;
  wire n6730_o;
  wire n6731_o;
  wire n6732_o;
  wire n6734_o;
  wire n6736_o;
  wire n6738_o;
  wire n6739_o;
  wire [5:0] n6740_o;
  wire n6742_o;
  wire [3:0] n6743_o;
  wire n6745_o;
  wire [1:0] n6746_o;
  wire n6748_o;
  wire n6749_o;
  wire n6750_o;
  wire n6755_o;
  wire n6758_o;
  wire n6761_o;
  wire n6764_o;
  wire n6765_o;
  wire n6766_o;
  wire n6768_o;
  wire n6769_o;
  wire n6770_o;
  wire n6771_o;
  wire n6772_o;
  wire n6773_o;
  wire n6774_o;
  wire n6775_o;
  wire n6776_o;
  wire n6777_o;
  wire n6778_o;
  wire n6779_o;
  wire n6780_o;
  wire [1:0] n6781_o;
  wire n6782_o;
  wire n6784_o;
  wire n6785_o;
  wire n6786_o;
  wire n6788_o;
  wire n6789_o;
  wire n6790_o;
  wire [1:0] n6791_o;
  wire n6793_o;
  wire n6795_o;
  wire n6797_o;
  wire n6799_o;
  wire n6800_o;
  wire n6801_o;
  wire n6802_o;
  wire n6804_o;
  wire n6805_o;
  wire n6806_o;
  wire n6807_o;
  wire n6808_o;
  wire n6809_o;
  wire n6810_o;
  wire n6811_o;
  wire [1:0] n6812_o;
  wire n6813_o;
  wire n6815_o;
  wire n6816_o;
  wire n6817_o;
  wire n6819_o;
  wire n6821_o;
  wire [6:0] n6822_o;
  wire n6824_o;
  wire [1:0] n6825_o;
  wire n6827_o;
  wire [2:0] n6828_o;
  wire n6830_o;
  wire n6832_o;
  wire [3:0] n6833_o;
  wire n6835_o;
  wire [1:0] n6836_o;
  wire n6838_o;
  wire n6839_o;
  wire n6840_o;
  wire [1:0] n6841_o;
  wire n6843_o;
  wire n6846_o;
  wire n6848_o;
  wire n6849_o;
  wire [1:0] n6850_o;
  wire n6852_o;
  wire n6853_o;
  wire n6854_o;
  wire n6858_o;
  wire n6860_o;
  wire [1:0] n6862_o;
  wire n6864_o;
  wire n6865_o;
  wire n6866_o;
  wire n6869_o;
  wire [1:0] n6872_o;
  wire [1:0] n6874_o;
  wire n6876_o;
  wire n6879_o;
  wire n6881_o;
  wire n6884_o;
  wire n6887_o;
  wire n6890_o;
  wire n6892_o;
  wire n6894_o;
  wire n6896_o;
  wire n6897_o;
  wire [1:0] n6898_o;
  wire n6900_o;
  wire n6901_o;
  wire [1:0] n6902_o;
  wire n6904_o;
  wire [3:0] n6907_o;
  wire n6909_o;
  wire [4:0] n6910_o;
  wire n6912_o;
  wire n6913_o;
  wire n6917_o;
  wire n6918_o;
  wire n6919_o;
  wire n6922_o;
  wire n6925_o;
  wire [1:0] n6927_o;
  wire n6930_o;
  wire [1:0] n6932_o;
  wire n6933_o;
  wire n6935_o;
  wire n6937_o;
  wire n6939_o;
  wire n6942_o;
  wire n6945_o;
  wire n6946_o;
  wire n6947_o;
  wire n6948_o;
  wire n6949_o;
  wire n6950_o;
  wire n6951_o;
  wire [1:0] n6952_o;
  wire [1:0] n6953_o;
  wire n6955_o;
  wire n6957_o;
  wire n6959_o;
  wire n6961_o;
  wire n6963_o;
  wire n6966_o;
  wire n6967_o;
  wire n6968_o;
  wire n6969_o;
  wire n6970_o;
  wire n6971_o;
  wire n6972_o;
  wire n6974_o;
  wire n6976_o;
  wire [1:0] n6977_o;
  wire n6979_o;
  wire n6980_o;
  wire n6981_o;
  wire [2:0] n6982_o;
  wire n6984_o;
  wire n6985_o;
  wire [3:0] n6986_o;
  wire n6988_o;
  wire [1:0] n6989_o;
  wire n6991_o;
  wire n6992_o;
  wire n6993_o;
  wire n6994_o;
  wire [1:0] n6995_o;
  wire n6997_o;
  wire n6998_o;
  wire [2:0] n6999_o;
  wire n7001_o;
  wire [1:0] n7002_o;
  wire n7004_o;
  wire n7005_o;
  wire n7006_o;
  wire n7007_o;
  wire n7008_o;
  wire n7012_o;
  wire n7015_o;
  wire n7018_o;
  wire n7020_o;
  wire [1:0] n7021_o;
  wire [1:0] n7022_o;
  wire n7024_o;
  wire n7026_o;
  wire n7028_o;
  wire n7029_o;
  wire n7030_o;
  wire n7032_o;
  wire n7034_o;
  wire n7035_o;
  wire n7036_o;
  wire n7037_o;
  wire n7038_o;
  wire n7039_o;
  wire n7040_o;
  wire n7042_o;
  wire n7044_o;
  wire n7046_o;
  wire [1:0] n7047_o;
  wire [1:0] n7048_o;
  wire n7050_o;
  wire n7052_o;
  wire n7054_o;
  wire n7056_o;
  wire n7057_o;
  wire n7058_o;
  wire n7059_o;
  wire n7061_o;
  wire n7063_o;
  wire n7065_o;
  wire n7066_o;
  wire n7067_o;
  wire n7068_o;
  wire n7069_o;
  wire n7070_o;
  wire n7071_o;
  wire n7073_o;
  wire n7075_o;
  wire n7077_o;
  wire n7079_o;
  wire n7081_o;
  wire n7083_o;
  wire n7085_o;
  wire [1:0] n7086_o;
  wire n7088_o;
  wire n7089_o;
  wire n7090_o;
  wire [1:0] n7091_o;
  wire n7093_o;
  wire [2:0] n7094_o;
  wire n7096_o;
  wire [1:0] n7097_o;
  wire n7099_o;
  wire n7100_o;
  wire n7101_o;
  wire [1:0] n7103_o;
  wire [1:0] n7106_o;
  wire n7109_o;
  wire [1:0] n7110_o;
  wire n7113_o;
  wire n7116_o;
  wire n7119_o;
  wire n7121_o;
  wire n7123_o;
  wire n7124_o;
  wire n7125_o;
  wire n7127_o;
  wire n7129_o;
  wire [1:0] n7130_o;
  wire n7132_o;
  wire [2:0] n7133_o;
  wire n7135_o;
  wire n7136_o;
  wire [2:0] n7137_o;
  wire n7139_o;
  wire n7140_o;
  wire [2:0] n7141_o;
  wire n7143_o;
  wire [2:0] n7144_o;
  wire n7146_o;
  wire n7147_o;
  wire [2:0] n7148_o;
  wire n7150_o;
  wire n7151_o;
  wire [2:0] n7152_o;
  wire n7154_o;
  wire [1:0] n7155_o;
  wire n7157_o;
  wire n7158_o;
  wire n7159_o;
  wire n7160_o;
  wire n7161_o;
  wire [1:0] n7162_o;
  wire n7164_o;
  wire [2:0] n7165_o;
  wire n7167_o;
  wire n7168_o;
  wire [2:0] n7169_o;
  wire n7171_o;
  wire n7172_o;
  wire [2:0] n7173_o;
  wire n7175_o;
  wire [2:0] n7176_o;
  wire n7178_o;
  wire n7179_o;
  wire [2:0] n7180_o;
  wire n7182_o;
  wire n7183_o;
  wire [3:0] n7184_o;
  wire n7186_o;
  wire n7187_o;
  wire n7188_o;
  wire n7189_o;
  wire n7192_o;
  wire n7193_o;
  wire n7194_o;
  wire n7195_o;
  wire [6:0] n7197_o;
  wire n7199_o;
  wire n7200_o;
  wire n7201_o;
  wire n7202_o;
  wire n7205_o;
  wire [2:0] n7206_o;
  wire n7208_o;
  wire n7211_o;
  wire [2:0] n7212_o;
  wire n7214_o;
  wire [2:0] n7215_o;
  wire n7217_o;
  wire n7218_o;
  wire [2:0] n7219_o;
  wire n7221_o;
  wire n7222_o;
  wire [2:0] n7223_o;
  wire n7225_o;
  wire n7226_o;
  wire n7229_o;
  wire [2:0] n7230_o;
  wire n7232_o;
  wire [2:0] n7233_o;
  wire n7235_o;
  wire n7236_o;
  wire [2:0] n7237_o;
  wire n7239_o;
  wire n7240_o;
  wire n7243_o;
  wire [1:0] n7244_o;
  wire n7246_o;
  wire [2:0] n7247_o;
  wire n7249_o;
  wire n7251_o;
  wire n7252_o;
  wire [1:0] n7255_o;
  wire n7258_o;
  wire n7261_o;
  wire n7262_o;
  wire n7263_o;
  wire n7264_o;
  wire n7266_o;
  wire n7268_o;
  wire n7270_o;
  wire n7271_o;
  wire n7272_o;
  wire [1:0] n7274_o;
  wire n7275_o;
  wire [1:0] n7279_o;
  wire n7281_o;
  wire n7283_o;
  wire n7284_o;
  wire n7285_o;
  wire n7286_o;
  wire [6:0] n7288_o;
  wire [2:0] n7289_o;
  wire n7291_o;
  wire n7294_o;
  wire n7297_o;
  wire [2:0] n7298_o;
  wire n7300_o;
  wire [2:0] n7301_o;
  wire n7303_o;
  wire n7304_o;
  wire [2:0] n7305_o;
  wire n7307_o;
  wire n7308_o;
  wire n7310_o;
  wire n7312_o;
  wire n7314_o;
  wire n7315_o;
  wire [1:0] n7316_o;
  wire n7318_o;
  wire n7321_o;
  wire n7323_o;
  wire n7325_o;
  wire n7327_o;
  wire n7329_o;
  wire n7332_o;
  wire n7335_o;
  wire n7336_o;
  wire n7337_o;
  wire n7338_o;
  wire n7339_o;
  wire n7340_o;
  wire n7341_o;
  wire n7342_o;
  wire n7343_o;
  wire [1:0] n7344_o;
  wire n7346_o;
  wire n7348_o;
  wire [1:0] n7350_o;
  wire [6:0] n7351_o;
  wire n7352_o;
  wire [1:0] n7353_o;
  wire n7354_o;
  wire n7356_o;
  wire n7358_o;
  wire n7360_o;
  wire n7362_o;
  wire n7364_o;
  wire n7365_o;
  wire n7366_o;
  wire n7367_o;
  wire n7369_o;
  wire n7370_o;
  wire n7371_o;
  wire n7372_o;
  wire n7373_o;
  wire n7374_o;
  wire n7375_o;
  wire n7376_o;
  wire n7377_o;
  wire n7378_o;
  wire n7380_o;
  wire [1:0] n7382_o;
  wire n7384_o;
  wire [6:0] n7385_o;
  wire n7391_o;
  wire [1:0] n7392_o;
  wire n7395_o;
  wire n7397_o;
  wire n7399_o;
  wire n7401_o;
  wire n7403_o;
  wire n7405_o;
  wire n7407_o;
  wire n7408_o;
  wire n7410_o;
  wire n7412_o;
  wire n7414_o;
  wire n7415_o;
  wire n7416_o;
  wire n7417_o;
  wire n7418_o;
  wire n7419_o;
  wire n7420_o;
  wire n7421_o;
  wire n7422_o;
  wire n7424_o;
  wire n7425_o;
  wire [1:0] n7427_o;
  wire n7428_o;
  wire [6:0] n7429_o;
  wire n7431_o;
  wire n7432_o;
  wire [2:0] n7433_o;
  wire n7435_o;
  wire n7436_o;
  wire [1:0] n7437_o;
  wire n7439_o;
  wire [2:0] n7440_o;
  wire n7442_o;
  wire n7443_o;
  wire [2:0] n7444_o;
  wire n7446_o;
  wire [1:0] n7447_o;
  wire n7449_o;
  wire n7450_o;
  wire n7451_o;
  wire [2:0] n7452_o;
  wire n7454_o;
  wire n7455_o;
  wire n7456_o;
  wire [1:0] n7457_o;
  wire n7459_o;
  wire n7460_o;
  wire n7463_o;
  wire n7466_o;
  wire n7468_o;
  wire n7471_o;
  wire n7473_o;
  wire n7476_o;
  wire n7479_o;
  wire n7481_o;
  wire n7482_o;
  wire n7483_o;
  wire n7485_o;
  wire n7487_o;
  wire n7489_o;
  wire n7490_o;
  wire [2:0] n7491_o;
  wire n7493_o;
  wire n7494_o;
  wire [1:0] n7495_o;
  wire n7497_o;
  wire [2:0] n7498_o;
  wire n7500_o;
  wire n7501_o;
  wire [2:0] n7502_o;
  wire n7504_o;
  wire [1:0] n7505_o;
  wire n7507_o;
  wire [2:0] n7508_o;
  wire n7510_o;
  wire n7511_o;
  wire n7512_o;
  wire n7513_o;
  wire [4:0] n7514_o;
  wire n7516_o;
  wire [2:0] n7517_o;
  wire n7519_o;
  wire [2:0] n7520_o;
  wire n7522_o;
  wire n7523_o;
  wire [2:0] n7524_o;
  wire n7526_o;
  wire n7529_o;
  wire n7532_o;
  wire n7534_o;
  wire n7537_o;
  wire n7539_o;
  wire n7542_o;
  wire n7545_o;
  wire n7547_o;
  wire n7548_o;
  wire n7549_o;
  wire n7551_o;
  wire n7553_o;
  wire n7555_o;
  wire n7557_o;
  wire n7559_o;
  wire n7561_o;
  wire n7563_o;
  wire n7565_o;
  wire n7567_o;
  wire n7568_o;
  wire n7569_o;
  wire n7570_o;
  wire n7572_o;
  wire [12:0] n7573_o;
  reg n7574_o;
  reg [1:0] n7576_o;
  reg [1:0] n7577_o;
  reg [1:0] n7578_o;
  reg n7579_o;
  reg n7581_o;
  reg n7582_o;
  reg n7584_o;
  reg n7586_o;
  reg n7587_o;
  reg n7589_o;
  reg n7591_o;
  reg n7593_o;
  reg n7595_o;
  reg n7597_o;
  reg n7599_o;
  reg n7601_o;
  reg n7603_o;
  reg n7605_o;
  reg n7607_o;
  reg [1:0] n7608_o;
  reg [5:0] n7609_o;
  reg n7611_o;
  reg n7612_o;
  reg n7615_o;
  reg n7617_o;
  reg n7620_o;
  reg n7622_o;
  reg n7624_o;
  reg n7626_o;
  reg n7631_o;
  reg n7633_o;
  reg n7635_o;
  reg n7637_o;
  reg n7639_o;
  reg n7641_o;
  wire n7642_o;
  reg n7643_o;
  wire [2:0] n7644_o;
  reg [2:0] n7645_o;
  wire n7646_o;
  reg n7647_o;
  wire n7648_o;
  reg n7649_o;
  wire n7650_o;
  reg n7651_o;
  wire n7652_o;
  reg n7653_o;
  wire n7654_o;
  reg n7655_o;
  wire n7656_o;
  reg n7657_o;
  wire n7658_o;
  reg n7659_o;
  reg n7660_o;
  wire n7661_o;
  reg n7662_o;
  wire n7663_o;
  reg n7664_o;
  wire n7665_o;
  wire n7666_o;
  reg n7667_o;
  wire n7668_o;
  wire n7669_o;
  reg n7670_o;
  wire n7671_o;
  reg n7672_o;
  wire n7673_o;
  wire n7674_o;
  wire n7675_o;
  wire n7676_o;
  wire n7677_o;
  reg n7678_o;
  wire n7679_o;
  wire n7680_o;
  wire n7681_o;
  wire n7682_o;
  wire n7683_o;
  reg n7684_o;
  wire n7685_o;
  wire n7686_o;
  reg n7687_o;
  wire n7688_o;
  wire n7689_o;
  reg n7690_o;
  wire n7691_o;
  reg n7692_o;
  wire [1:0] n7693_o;
  wire [1:0] n7694_o;
  reg [1:0] n7695_o;
  wire n7696_o;
  wire n7697_o;
  reg n7698_o;
  wire n7699_o;
  wire n7700_o;
  reg n7701_o;
  wire n7702_o;
  wire n7703_o;
  wire n7704_o;
  reg n7705_o;
  wire n7706_o;
  wire n7707_o;
  reg n7708_o;
  wire [3:0] n7709_o;
  reg [3:0] n7710_o;
  wire n7711_o;
  reg n7712_o;
  wire n7713_o;
  wire [4:0] n7714_o;
  reg [4:0] n7715_o;
  wire n7716_o;
  reg n7717_o;
  wire n7718_o;
  reg n7719_o;
  wire n7720_o;
  reg n7721_o;
  wire n7722_o;
  wire n7723_o;
  reg n7724_o;
  wire n7725_o;
  reg n7726_o;
  wire n7727_o;
  reg n7728_o;
  wire n7729_o;
  reg n7730_o;
  wire n7731_o;
  reg n7732_o;
  wire n7733_o;
  reg n7734_o;
  wire n7735_o;
  reg n7737_o;
  wire n7738_o;
  reg n7740_o;
  wire n7741_o;
  reg n7743_o;
  wire n7744_o;
  wire n7745_o;
  reg n7747_o;
  wire n7748_o;
  reg n7750_o;
  wire n7751_o;
  reg n7753_o;
  wire n7754_o;
  wire n7755_o;
  reg n7757_o;
  wire n7758_o;
  wire n7759_o;
  reg n7761_o;
  wire n7762_o;
  reg n7764_o;
  reg n7766_o;
  reg n7768_o;
  reg n7770_o;
  reg n7772_o;
  reg n7774_o;
  reg n7776_o;
  reg n7778_o;
  reg n7780_o;
  reg n7782_o;
  reg n7784_o;
  reg n7786_o;
  reg n7788_o;
  reg [1:0] n7790_o;
  reg n7792_o;
  reg n7794_o;
  reg [1:0] n7796_o;
  reg [1:0] n7798_o;
  reg n7800_o;
  reg n7802_o;
  reg [6:0] n7803_o;
  wire n7804_o;
  wire [1:0] n7805_o;
  wire [1:0] n7806_o;
  wire [1:0] n7807_o;
  wire n7808_o;
  wire n7810_o;
  wire n7812_o;
  wire n7814_o;
  wire n7817_o;
  wire n7819_o;
  wire n7821_o;
  wire n7824_o;
  wire n7827_o;
  wire n7830_o;
  wire n7833_o;
  wire n7836_o;
  wire n7839_o;
  wire n7842_o;
  wire n7845_o;
  wire n7848_o;
  wire [1:0] n7850_o;
  wire [5:0] n7851_o;
  wire n7853_o;
  wire n7855_o;
  wire n7857_o;
  wire n7861_o;
  wire n7864_o;
  wire n7867_o;
  wire n7870_o;
  wire n7873_o;
  wire n7876_o;
  wire n7879_o;
  wire n7882_o;
  wire n7885_o;
  wire n7888_o;
  wire n7891_o;
  wire n7894_o;
  wire [3:0] n7896_o;
  wire [4:0] n7897_o;
  wire [2:0] n7898_o;
  wire [15:0] n7899_o;
  wire [1:0] n7900_o;
  wire [2:0] n7901_o;
  wire n7902_o;
  wire n7903_o;
  wire n7906_o;
  wire n7907_o;
  wire n7908_o;
  wire n7909_o;
  wire n7910_o;
  wire n7911_o;
  wire n7912_o;
  wire n7913_o;
  wire [1:0] n7914_o;
  wire [4:0] n7915_o;
  wire [2:0] n7917_o;
  wire [2:0] n7918_o;
  wire [15:0] n7919_o;
  wire n7921_o;
  wire [4:0] n7922_o;
  wire n7924_o;
  wire n7925_o;
  wire n7926_o;
  wire n7927_o;
  wire n7928_o;
  wire [1:0] n7929_o;
  wire n7931_o;
  wire n7932_o;
  wire n7933_o;
  wire n7934_o;
  wire n7938_o;
  wire [15:0] n7939_o;
  wire n7940_o;
  wire [3:0] n7945_o;
  wire n7946_o;
  wire n7947_o;
  wire n7950_o;
  wire n7951_o;
  wire n7952_o;
  wire n7956_o;
  wire [8:0] n7958_o;
  wire [6:0] n7959_o;
  wire [4:0] n7960_o;
  wire [3:0] n7961_o;
  wire [8:0] n7963_o;
  wire [6:0] n7965_o;
  wire n7967_o;
  wire n7969_o;
  wire n7971_o;
  localparam [4:0] n7972_o = 5'b00000;
  wire n7975_o;
  wire [3:0] n7977_o;
  wire n7979_o;
  wire n7981_o;
  localparam [88:0] n7982_o = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n7985_o;
  wire [2:0] n7987_o;
  wire n7991_o;
  wire n7993_o;
  wire [31:0] n7995_o;
  wire [6:0] n7997_o;
  wire [1:0] n7999_o;
  wire [5:0] n8000_o;
  wire [6:0] n8001_o;
  wire n8002_o;
  wire n8003_o;
  wire n8004_o;
  wire n8005_o;
  wire [1:0] n8006_o;
  wire n8008_o;
  wire n8009_o;
  wire n8010_o;
  wire n8012_o;
  wire n8013_o;
  wire n8014_o;
  wire n8015_o;
  wire n8016_o;
  wire n8018_o;
  wire n8020_o;
  wire n8022_o;
  wire n8024_o;
  wire n8025_o;
  wire n8027_o;
  wire n8028_o;
  wire n8029_o;
  wire n8030_o;
  wire n8031_o;
  wire n8032_o;
  wire n8033_o;
  wire n8035_o;
  wire n8036_o;
  wire n8037_o;
  wire n8038_o;
  wire n8039_o;
  wire n8040_o;
  wire [3:0] n8041_o;
  wire [3:0] n8042_o;
  wire [3:0] n8043_o;
  wire n8046_o;
  wire [2:0] n8047_o;
  wire n8049_o;
  wire n8051_o;
  wire n8052_o;
  wire n8053_o;
  wire n8054_o;
  wire [1:0] n8058_o;
  wire n8060_o;
  wire n8061_o;
  wire n8062_o;
  wire n8063_o;
  wire n8064_o;
  wire n8065_o;
  wire n8066_o;
  wire n8067_o;
  wire n8068_o;
  wire n8069_o;
  wire n8070_o;
  wire n8071_o;
  wire n8072_o;
  wire [6:0] n8074_o;
  wire n8076_o;
  wire n8077_o;
  wire n8079_o;
  wire n8080_o;
  wire n8081_o;
  wire n8082_o;
  wire n8083_o;
  wire n8084_o;
  wire n8085_o;
  wire n8086_o;
  wire n8087_o;
  wire n8088_o;
  wire n8089_o;
  wire n8090_o;
  wire n8091_o;
  wire n8092_o;
  wire n8093_o;
  wire n8094_o;
  wire n8096_o;
  wire n8098_o;
  wire n8099_o;
  wire n8100_o;
  wire n8101_o;
  wire n8102_o;
  wire n8103_o;
  wire n8104_o;
  wire n8105_o;
  wire n8106_o;
  wire n8107_o;
  wire n8108_o;
  wire n8109_o;
  wire n8110_o;
  wire n8111_o;
  wire n8112_o;
  wire n8122_o;
  wire n8123_o;
  wire n8124_o;
  wire n8131_o;
  wire n8132_o;
  wire n8133_o;
  wire n8134_o;
  wire n8135_o;
  wire n8137_o;
  wire n8138_o;
  wire n8140_o;
  wire n8142_o;
  wire [6:0] n8143_o;
  wire n8144_o;
  wire [6:0] n8146_o;
  wire n8152_o;
  wire n8155_o;
  wire n8158_o;
  wire n8159_o;
  wire n8160_o;
  wire n8162_o;
  wire n8163_o;
  wire n8164_o;
  wire n8166_o;
  wire n8167_o;
  wire n8169_o;
  wire n8170_o;
  wire n8172_o;
  wire n8174_o;
  wire n8175_o;
  wire n8176_o;
  wire n8177_o;
  wire n8178_o;
  wire n8180_o;
  wire n8181_o;
  wire n8182_o;
  wire n8183_o;
  wire [1:0] n8185_o;
  wire n8186_o;
  wire n8187_o;
  wire n8188_o;
  wire n8189_o;
  wire [1:0] n8191_o;
  wire n8194_o;
  wire n8197_o;
  wire n8198_o;
  wire n8199_o;
  wire n8200_o;
  wire n8201_o;
  wire n8202_o;
  wire n8203_o;
  wire n8204_o;
  wire [6:0] n8207_o;
  wire n8209_o;
  wire n8212_o;
  wire n8213_o;
  wire n8216_o;
  wire n8217_o;
  wire n8218_o;
  wire n8219_o;
  wire n8220_o;
  wire n8221_o;
  wire [1:0] n8223_o;
  wire n8225_o;
  wire [6:0] n8228_o;
  wire [1:0] n8229_o;
  wire n8231_o;
  wire [1:0] n8235_o;
  wire n8238_o;
  wire n8240_o;
  wire n8241_o;
  wire n8242_o;
  wire n8243_o;
  wire n8244_o;
  wire n8245_o;
  wire [6:0] n8247_o;
  wire [1:0] n8249_o;
  wire n8251_o;
  wire n8252_o;
  wire n8253_o;
  wire n8254_o;
  wire n8255_o;
  wire n8256_o;
  wire n8257_o;
  wire n8258_o;
  wire [6:0] n8259_o;
  wire n8261_o;
  wire n8264_o;
  wire n8266_o;
  wire n8267_o;
  wire n8268_o;
  wire n8270_o;
  wire n8271_o;
  wire n8272_o;
  wire n8273_o;
  wire [1:0] n8275_o;
  wire n8276_o;
  wire n8277_o;
  wire n8278_o;
  wire n8279_o;
  wire n8281_o;
  wire n8282_o;
  wire n8285_o;
  wire n8286_o;
  wire n8287_o;
  wire n8288_o;
  wire n8289_o;
  wire [1:0] n8293_o;
  wire n8295_o;
  wire n8296_o;
  wire n8297_o;
  wire [6:0] n8299_o;
  wire n8301_o;
  wire n8303_o;
  wire n8304_o;
  wire n8305_o;
  wire n8307_o;
  wire n8308_o;
  wire n8309_o;
  wire n8311_o;
  wire n8312_o;
  wire n8314_o;
  wire n8316_o;
  wire n8317_o;
  wire n8318_o;
  wire n8319_o;
  wire n8321_o;
  wire n8322_o;
  wire n8323_o;
  wire n8324_o;
  wire [1:0] n8326_o;
  wire n8327_o;
  wire n8328_o;
  wire n8329_o;
  wire n8330_o;
  wire [1:0] n8332_o;
  wire n8335_o;
  wire n8338_o;
  wire n8339_o;
  wire n8340_o;
  wire n8341_o;
  wire n8342_o;
  wire n8343_o;
  wire n8344_o;
  wire [6:0] n8347_o;
  wire n8349_o;
  wire n8352_o;
  wire n8353_o;
  wire n8356_o;
  wire n8357_o;
  wire n8358_o;
  wire n8359_o;
  wire n8360_o;
  wire n8361_o;
  wire [1:0] n8363_o;
  wire n8365_o;
  wire [6:0] n8368_o;
  wire [1:0] n8369_o;
  wire n8371_o;
  wire [1:0] n8376_o;
  wire n8377_o;
  wire n8378_o;
  wire n8379_o;
  wire n8380_o;
  wire n8381_o;
  wire n8382_o;
  wire n8383_o;
  wire n8384_o;
  wire [6:0] n8387_o;
  wire [1:0] n8389_o;
  wire n8390_o;
  wire n8391_o;
  wire n8392_o;
  wire n8393_o;
  wire n8394_o;
  wire n8395_o;
  wire n8396_o;
  wire n8397_o;
  wire n8398_o;
  wire [6:0] n8399_o;
  wire n8401_o;
  wire n8405_o;
  wire n8408_o;
  wire n8409_o;
  wire n8410_o;
  wire n8412_o;
  wire n8413_o;
  wire n8414_o;
  wire n8415_o;
  wire [1:0] n8417_o;
  wire n8418_o;
  wire n8419_o;
  wire n8420_o;
  wire n8421_o;
  wire n8423_o;
  wire n8425_o;
  wire n8428_o;
  wire n8429_o;
  wire n8430_o;
  wire n8431_o;
  wire n8432_o;
  wire [1:0] n8436_o;
  wire n8437_o;
  wire [6:0] n8440_o;
  wire n8442_o;
  wire n8444_o;
  wire n8447_o;
  wire [6:0] n8449_o;
  wire n8451_o;
  wire n8453_o;
  wire n8454_o;
  wire n8457_o;
  wire n8460_o;
  wire n8462_o;
  wire n8463_o;
  wire n8464_o;
  wire n8466_o;
  wire n8469_o;
  wire [6:0] n8471_o;
  wire n8472_o;
  wire n8475_o;
  wire n8477_o;
  wire n8478_o;
  wire n8480_o;
  wire n8486_o;
  wire n8487_o;
  wire [1:0] n8488_o;
  wire n8490_o;
  wire n8492_o;
  wire n8493_o;
  wire [1:0] n8495_o;
  wire n8498_o;
  wire n8500_o;
  wire n8505_o;
  wire n8507_o;
  wire [1:0] n8509_o;
  wire n8512_o;
  wire n8516_o;
  wire n8517_o;
  wire [1:0] n8519_o;
  wire [6:0] n8521_o;
  wire n8523_o;
  wire n8525_o;
  wire n8526_o;
  wire n8528_o;
  wire n8530_o;
  wire n8532_o;
  wire n8533_o;
  wire [1:0] n8540_o;
  wire n8543_o;
  wire n8544_o;
  wire n8545_o;
  wire n8546_o;
  wire n8547_o;
  wire n8548_o;
  wire n8549_o;
  wire n8550_o;
  wire n8551_o;
  wire n8552_o;
  wire n8553_o;
  wire n8554_o;
  wire n8555_o;
  wire [6:0] n8557_o;
  wire n8559_o;
  wire n8560_o;
  wire n8563_o;
  wire n8569_o;
  wire n8572_o;
  wire n8573_o;
  wire n8575_o;
  wire n8576_o;
  wire n8577_o;
  wire n8578_o;
  wire n8584_o;
  wire n8587_o;
  wire n8588_o;
  wire n8590_o;
  wire [1:0] n8598_o;
  wire n8601_o;
  wire n8603_o;
  wire n8606_o;
  wire n8608_o;
  wire n8609_o;
  wire n8610_o;
  wire n8611_o;
  wire n8612_o;
  wire n8613_o;
  wire n8614_o;
  wire n8615_o;
  wire n8616_o;
  wire n8617_o;
  wire n8618_o;
  wire n8619_o;
  wire n8620_o;
  wire n8621_o;
  wire n8622_o;
  wire n8623_o;
  wire n8624_o;
  wire n8625_o;
  wire [6:0] n8628_o;
  wire n8630_o;
  wire n8634_o;
  wire n8638_o;
  wire [15:0] n8639_o;
  wire n8641_o;
  wire [2:0] n8642_o;
  wire n8644_o;
  wire n8646_o;
  wire n8648_o;
  wire n8649_o;
  wire n8650_o;
  wire n8651_o;
  wire n8652_o;
  wire n8653_o;
  wire [1:0] n8655_o;
  wire n8656_o;
  wire n8657_o;
  wire n8658_o;
  wire n8659_o;
  wire n8660_o;
  wire [6:0] n8662_o;
  wire n8664_o;
  wire n8665_o;
  wire n8668_o;
  wire n8669_o;
  wire [1:0] n8673_o;
  wire n8674_o;
  wire n8675_o;
  wire n8676_o;
  wire n8677_o;
  wire [1:0] n8679_o;
  wire n8680_o;
  wire n8681_o;
  wire n8682_o;
  wire n8683_o;
  wire n8684_o;
  wire n8685_o;
  wire n8686_o;
  wire n8687_o;
  wire n8688_o;
  wire [6:0] n8690_o;
  wire n8692_o;
  wire [1:0] n8693_o;
  wire n8695_o;
  wire n8697_o;
  wire n8699_o;
  wire [2:0] n8700_o;
  wire n8702_o;
  wire n8704_o;
  wire n8709_o;
  wire [2:0] n8710_o;
  wire n8712_o;
  wire n8714_o;
  wire [1:0] n8716_o;
  wire n8718_o;
  wire [1:0] n8721_o;
  wire n8724_o;
  wire n8726_o;
  wire [2:0] n8727_o;
  wire n8729_o;
  wire n8731_o;
  wire n8734_o;
  wire [2:0] n8735_o;
  wire n8737_o;
  wire n8739_o;
  wire n8742_o;
  wire n8746_o;
  wire n8749_o;
  wire n8752_o;
  wire n8755_o;
  wire n8758_o;
  wire n8761_o;
  wire n8762_o;
  wire n8764_o;
  wire [1:0] n8767_o;
  wire n8768_o;
  wire n8769_o;
  wire [6:0] n8772_o;
  wire n8774_o;
  wire n8775_o;
  wire n8777_o;
  wire n8780_o;
  wire n8783_o;
  wire n8787_o;
  wire n8790_o;
  wire n8793_o;
  wire n8796_o;
  wire n8799_o;
  wire n8802_o;
  wire n8805_o;
  wire n8808_o;
  wire n8811_o;
  wire n8812_o;
  wire n8813_o;
  wire n8816_o;
  wire n8817_o;
  wire n8818_o;
  wire n8819_o;
  wire n8820_o;
  wire n8822_o;
  wire n8824_o;
  wire n8825_o;
  wire n8826_o;
  wire [1:0] n8829_o;
  wire n8831_o;
  wire n8832_o;
  wire [6:0] n8835_o;
  wire n8837_o;
  wire n8839_o;
  wire [3:0] n8840_o;
  wire n8842_o;
  wire [1:0] n8846_o;
  wire [1:0] n8848_o;
  wire n8850_o;
  wire n8851_o;
  wire [6:0] n8854_o;
  wire n8856_o;
  wire n8858_o;
  wire n8860_o;
  wire n8863_o;
  wire [11:0] n8865_o;
  wire n8867_o;
  wire [11:0] n8868_o;
  wire n8870_o;
  wire n8871_o;
  wire [11:0] n8872_o;
  wire n8874_o;
  wire n8875_o;
  wire [11:0] n8876_o;
  wire n8878_o;
  wire n8879_o;
  wire n8880_o;
  wire [11:0] n8881_o;
  wire n8883_o;
  wire [11:0] n8884_o;
  wire n8886_o;
  wire n8887_o;
  wire [11:0] n8888_o;
  wire n8890_o;
  wire n8891_o;
  wire [11:0] n8892_o;
  wire n8894_o;
  wire n8895_o;
  wire n8896_o;
  wire n8897_o;
  wire n8898_o;
  wire n8899_o;
  wire n8901_o;
  wire n8903_o;
  wire n8905_o;
  wire n8906_o;
  wire n8908_o;
  wire n8912_o;
  wire n8914_o;
  wire n8915_o;
  wire n8916_o;
  wire n8917_o;
  wire n8918_o;
  wire n8919_o;
  wire [1:0] n8922_o;
  wire n8924_o;
  wire n8925_o;
  wire n8928_o;
  wire n8929_o;
  wire n8930_o;
  wire n8931_o;
  wire n8932_o;
  wire n8933_o;
  wire n8934_o;
  wire n8935_o;
  wire n8936_o;
  wire n8937_o;
  wire [1:0] n8940_o;
  wire n8942_o;
  wire n8943_o;
  wire n8947_o;
  wire n8948_o;
  wire [1:0] n8951_o;
  wire [1:0] n8953_o;
  wire [1:0] n8954_o;
  wire n8955_o;
  wire n8956_o;
  wire n8957_o;
  wire n8958_o;
  wire n8959_o;
  wire n8960_o;
  wire n8961_o;
  wire n8962_o;
  wire n8963_o;
  wire [6:0] n8965_o;
  wire n8967_o;
  wire n8968_o;
  wire n8969_o;
  wire [1:0] n8972_o;
  wire n8974_o;
  wire n8976_o;
  wire n8977_o;
  wire n8979_o;
  wire [5:0] n8982_o;
  wire n8984_o;
  wire n8987_o;
  wire [6:0] n8990_o;
  wire n8992_o;
  wire n8993_o;
  wire n8994_o;
  wire n8996_o;
  wire n8998_o;
  wire n8999_o;
  wire n9001_o;
  wire n9003_o;
  wire [1:0] n9005_o;
  wire [6:0] n9007_o;
  wire n9009_o;
  wire n9011_o;
  wire n9012_o;
  wire n9013_o;
  wire n9014_o;
  wire n9015_o;
  wire n9016_o;
  wire n9017_o;
  wire n9019_o;
  wire n9024_o;
  wire n9026_o;
  wire [15:0] n9027_o;
  wire n9029_o;
  wire n9030_o;
  wire n9031_o;
  wire n9033_o;
  wire [15:0] n9034_o;
  wire n9036_o;
  wire n9037_o;
  wire n9040_o;
  wire [6:0] n9042_o;
  wire n9045_o;
  wire n9046_o;
  wire n9048_o;
  wire [5:0] n9051_o;
  wire n9053_o;
  wire n9056_o;
  wire [6:0] n9059_o;
  wire n9061_o;
  wire n9062_o;
  wire n9063_o;
  wire n9064_o;
  wire n9066_o;
  wire n9067_o;
  wire n9068_o;
  wire n9070_o;
  wire [1:0] n9073_o;
  wire n9076_o;
  wire n9077_o;
  wire [6:0] n9079_o;
  wire n9082_o;
  wire n9083_o;
  wire n9086_o;
  wire n9087_o;
  wire n9088_o;
  wire n9089_o;
  wire n9090_o;
  wire n9093_o;
  wire [5:0] n9094_o;
  wire n9096_o;
  wire [5:0] n9097_o;
  wire [5:0] n9099_o;
  wire n9100_o;
  wire n9101_o;
  wire n9103_o;
  wire n9105_o;
  wire [84:0] n9106_o;
  reg n9109_o;
  reg [1:0] n9126_o;
  reg [1:0] n9127_o;
  reg [1:0] n9169_o;
  reg n9172_o;
  reg n9175_o;
  reg n9180_o;
  reg n9182_o;
  reg n9192_o;
  reg n9196_o;
  reg n9214_o;
  reg n9216_o;
  reg n9219_o;
  reg n9222_o;
  reg n9225_o;
  reg n9229_o;
  reg n9233_o;
  reg n9236_o;
  reg n9241_o;
  reg n9243_o;
  reg n9248_o;
  reg n9251_o;
  reg n9257_o;
  reg n9261_o;
  reg n9266_o;
  reg [5:0] n9267_o;
  reg n9271_o;
  reg n9274_o;
  reg n9278_o;
  reg n9280_o;
  reg n9281_o;
  reg n9284_o;
  reg n9286_o;
  reg n9288_o;
  wire n9289_o;
  wire n9290_o;
  wire n9291_o;
  reg n9292_o;
  reg n9293_o;
  reg n9294_o;
  reg n9295_o;
  reg n9296_o;
  reg n9297_o;
  wire n9298_o;
  reg n9299_o;
  reg n9300_o;
  reg n9301_o;
  wire n9302_o;
  wire n9303_o;
  wire n9304_o;
  reg n9305_o;
  reg n9306_o;
  wire n9307_o;
  wire n9308_o;
  wire n9309_o;
  reg n9310_o;
  wire n9311_o;
  wire n9312_o;
  wire n9313_o;
  reg n9314_o;
  reg n9315_o;
  reg n9316_o;
  reg n9317_o;
  wire n9318_o;
  wire n9319_o;
  wire n9320_o;
  reg n9321_o;
  reg n9322_o;
  wire n9323_o;
  wire n9324_o;
  wire n9325_o;
  reg n9326_o;
  wire n9327_o;
  wire n9328_o;
  wire n9329_o;
  reg n9330_o;
  wire n9331_o;
  wire n9332_o;
  wire n9333_o;
  reg n9334_o;
  wire n9335_o;
  wire n9336_o;
  wire n9337_o;
  reg n9338_o;
  reg n9339_o;
  wire n9340_o;
  wire n9341_o;
  wire n9342_o;
  reg n9343_o;
  wire n9344_o;
  wire n9345_o;
  wire n9346_o;
  reg n9347_o;
  reg n9348_o;
  reg n9349_o;
  reg n9350_o;
  reg n9351_o;
  wire n9352_o;
  wire n9353_o;
  wire n9354_o;
  reg n9355_o;
  wire n9356_o;
  reg n9357_o;
  reg n9358_o;
  reg n9359_o;
  wire n9360_o;
  wire n9361_o;
  wire n9362_o;
  reg n9363_o;
  wire n9364_o;
  wire n9365_o;
  wire n9366_o;
  reg n9367_o;
  wire n9368_o;
  wire n9369_o;
  wire n9370_o;
  reg n9371_o;
  wire n9372_o;
  reg n9373_o;
  wire n9374_o;
  reg n9375_o;
  wire [2:0] n9376_o;
  wire [2:0] n9377_o;
  wire [2:0] n9378_o;
  wire n9379_o;
  wire n9380_o;
  wire n9381_o;
  wire n9382_o;
  wire n9386_o;
  wire n9387_o;
  wire n9388_o;
  wire [3:0] n9392_o;
  wire [3:0] n9393_o;
  wire [3:0] n9394_o;
  wire [2:0] n9401_o;
  wire [2:0] n9402_o;
  wire [2:0] n9403_o;
  wire n9407_o;
  wire n9408_o;
  wire n9409_o;
  wire [1:0] n9410_o;
  wire [1:0] n9411_o;
  wire [1:0] n9412_o;
  wire n9413_o;
  wire n9414_o;
  wire n9415_o;
  wire [3:0] n9416_o;
  wire n9424_o;
  reg n9425_o;
  wire [1:0] n9426_o;
  wire [1:0] n9427_o;
  reg [6:0] n9473_o;
  wire n9478_o;
  wire n9479_o;
  wire [11:0] n9480_o;
  wire [2:0] n9481_o;
  wire n9483_o;
  wire [2:0] n9484_o;
  wire n9486_o;
  wire [3:0] n9487_o;
  wire n9489_o;
  wire n9491_o;
  wire n9493_o;
  wire n9495_o;
  wire n9497_o;
  wire n9499_o;
  wire [7:0] n9500_o;
  reg [31:0] n9501_o;
  reg [3:0] n9502_o;
  reg [2:0] n9503_o;
  reg [2:0] n9504_o;
  wire [31:0] n9505_o;
  wire [3:0] n9506_o;
  wire [2:0] n9507_o;
  wire [2:0] n9508_o;
  wire [31:0] n9510_o;
  wire [3:0] n9512_o;
  wire [2:0] n9513_o;
  wire [2:0] n9514_o;
  wire [11:0] n9519_o;
  wire [31:0] n9521_o;
  wire n9523_o;
  wire [31:0] n9525_o;
  wire n9527_o;
  wire [3:0] n9529_o;
  wire [31:0] n9531_o;
  wire n9533_o;
  wire n9535_o;
  wire [3:0] n9536_o;
  reg [31:0] n9538_o;
  wire [3:0] n9543_o;
  wire n9545_o;
  wire n9547_o;
  wire n9548_o;
  wire n9549_o;
  wire n9550_o;
  wire n9551_o;
  wire n9552_o;
  wire n9554_o;
  wire n9555_o;
  wire n9556_o;
  wire n9557_o;
  wire n9559_o;
  wire n9560_o;
  wire n9561_o;
  wire n9563_o;
  wire n9564_o;
  wire n9566_o;
  wire n9567_o;
  wire n9568_o;
  wire n9570_o;
  wire n9571_o;
  wire n9573_o;
  wire n9574_o;
  wire n9575_o;
  wire n9577_o;
  wire n9578_o;
  wire n9580_o;
  wire n9581_o;
  wire n9582_o;
  wire n9584_o;
  wire n9585_o;
  wire n9587_o;
  wire n9588_o;
  wire n9589_o;
  wire n9590_o;
  wire n9591_o;
  wire n9592_o;
  wire n9593_o;
  wire n9594_o;
  wire n9595_o;
  wire n9596_o;
  wire n9598_o;
  wire n9599_o;
  wire n9600_o;
  wire n9601_o;
  wire n9602_o;
  wire n9603_o;
  wire n9604_o;
  wire n9605_o;
  wire n9606_o;
  wire n9607_o;
  wire n9609_o;
  wire n9610_o;
  wire n9611_o;
  wire n9612_o;
  wire n9613_o;
  wire n9614_o;
  wire n9615_o;
  wire n9616_o;
  wire n9617_o;
  wire n9618_o;
  wire n9619_o;
  wire n9620_o;
  wire n9621_o;
  wire n9622_o;
  wire n9623_o;
  wire n9624_o;
  wire n9626_o;
  wire n9627_o;
  wire n9628_o;
  wire n9629_o;
  wire n9630_o;
  wire n9631_o;
  wire n9632_o;
  wire n9633_o;
  wire n9634_o;
  wire n9635_o;
  wire n9636_o;
  wire n9637_o;
  wire n9639_o;
  wire [15:0] n9640_o;
  reg n9643_o;
  wire n9648_o;
  wire [15:0] n9649_o;
  wire n9650_o;
  wire n9651_o;
  wire n9652_o;
  wire n9655_o;
  wire n9658_o;
  wire n9661_o;
  wire n9664_o;
  wire n9667_o;
  wire n9670_o;
  wire n9673_o;
  wire n9676_o;
  wire n9679_o;
  wire n9682_o;
  wire n9685_o;
  wire n9688_o;
  wire n9691_o;
  wire n9694_o;
  wire n9697_o;
  wire n9700_o;
  wire [15:0] n9701_o;
  wire n9702_o;
  reg n9703_o;
  wire n9704_o;
  reg n9705_o;
  wire n9706_o;
  reg n9707_o;
  wire n9708_o;
  reg n9709_o;
  wire n9710_o;
  reg n9711_o;
  wire n9712_o;
  reg n9713_o;
  wire n9714_o;
  reg n9715_o;
  wire n9716_o;
  reg n9717_o;
  wire n9718_o;
  reg n9719_o;
  wire n9720_o;
  reg n9721_o;
  wire n9722_o;
  reg n9723_o;
  wire n9724_o;
  reg n9725_o;
  wire n9726_o;
  reg n9727_o;
  wire n9728_o;
  reg n9729_o;
  wire n9730_o;
  reg n9731_o;
  wire n9732_o;
  reg n9733_o;
  wire [15:0] n9734_o;
  wire [15:0] n9735_o;
  wire [15:0] n9736_o;
  wire [3:0] n9744_o;
  wire n9746_o;
  wire [3:0] n9747_o;
  wire n9749_o;
  wire [3:0] n9751_o;
  wire n9753_o;
  wire [3:0] n9754_o;
  wire n9756_o;
  wire n9759_o;
  wire [3:0] n9761_o;
  wire [3:0] n9762_o;
  wire n9764_o;
  wire [3:0] n9765_o;
  wire n9767_o;
  wire [3:0] n9768_o;
  wire [1:0] n9770_o;
  wire n9771_o;
  wire n9772_o;
  wire n9773_o;
  wire n9775_o;
  wire [3:0] n9776_o;
  wire n9778_o;
  wire [3:0] n9779_o;
  wire [1:0] n9780_o;
  wire [1:0] n9782_o;
  localparam [3:0] n9783_o = 4'b0000;
  wire [3:0] n9785_o;
  wire n9787_o;
  wire [1:0] n9789_o;
  wire n9791_o;
  wire n9793_o;
  wire n9794_o;
  wire n9796_o;
  wire n9797_o;
  wire n9798_o;
  wire n9799_o;
  wire n9801_o;
  wire n9802_o;
  wire [1:0] n9803_o;
  wire n9804_o;
  wire n9805_o;
  wire n9806_o;
  wire n9807_o;
  wire n9808_o;
  reg n9811_q;
  wire [3:0] n9812_o;
  reg [3:0] n9813_q;
  wire n9814_o;
  reg n9815_q;
  reg [31:0] n9816_q;
  wire [31:0] n9817_o;
  reg [31:0] n9818_q;
  wire [31:0] n9819_o;
  reg [31:0] n9820_q;
  reg [1:0] n9821_q;
  reg [1:0] n9822_q;
  reg n9823_q;
  reg [15:0] n9824_q;
  reg [15:0] n9825_q;
  wire [15:0] n9826_o;
  reg [15:0] n9827_q;
  reg [31:0] n9828_q;
  reg [31:0] n9829_q;
  reg [15:0] n9830_q;
  wire [3:0] n9832_o;
  reg [3:0] n9833_q;
  wire [31:0] n9834_o;
  wire [3:0] n9837_o;
  reg [3:0] n9838_q;
  wire [3:0] n9839_o;
  reg [3:0] n9840_q;
  wire n9841_o;
  reg n9842_q;
  wire [31:0] n9843_o;
  reg [31:0] n9844_q;
  wire [31:0] n9845_o;
  reg [31:0] n9846_q;
  wire n9847_o;
  reg n9848_q;
  reg [31:0] n9849_q;
  wire [31:0] n9850_o;
  reg [31:0] n9852_q;
  reg n9853_q;
  wire [31:0] n9855_o;
  reg n9856_q;
  reg [15:0] n9857_q;
  reg n9858_q;
  reg n9859_q;
  reg n9860_q;
  reg n9861_q;
  reg n9862_q;
  reg n9863_q;
  reg n9864_q;
  reg [7:0] n9865_q;
  reg n9866_q;
  wire n9867_o;
  reg n9868_q;
  reg [1:0] n9869_q;
  reg [5:0] n9870_q;
  wire n9871_o;
  reg n9872_q;
  wire [3:0] n9873_o;
  reg n9875_q;
  reg n9876_q;
  reg n9877_q;
  reg n9878_q;
  reg n9879_q;
  reg n9880_q;
  reg [7:0] n9881_q;
  reg n9882_q;
  reg n9883_q;
  reg n9884_q;
  reg n9885_q;
  wire [31:0] n9886_o;
  reg [31:0] n9887_q;
  wire [31:0] n9888_o;
  reg [31:0] n9889_q;
  reg [2:0] n9890_q;
  reg [7:0] n9891_q;
  reg n9892_q;
  reg n9893_q;
  reg n9894_q;
  reg n9895_q;
  reg n9896_q;
  wire [31:0] n9897_o;
  wire [7:0] n9898_o;
  reg [7:0] n9899_q;
  reg [5:0] n9900_q;
  reg [3:0] n9901_q;
  reg [5:0] n9902_q;
  reg n9903_q;
  reg n9904_q;
  reg [31:0] n9905_q;
  reg [31:0] n9906_q;
  wire [5:0] n9907_o;
  wire [5:0] n9908_o;
  reg [5:0] n9909_q;
  reg [5:0] n9910_q;
  wire [5:0] n9911_o;
  reg [31:0] n9912_q;
  reg [5:0] n9913_q;
  reg [31:0] n9914_q;
  reg [3:0] n9915_q;
  reg [2:0] n9916_q;
  reg [2:0] n9917_q;
  wire [88:0] n9918_o;
  wire [88:0] n9919_o;
  wire [88:0] n9920_o;
  reg [88:0] n9921_q;
  reg [6:0] n9922_q;
  reg n9923_q;
  reg [1:0] n9924_q;
  wire [2:0] n9925_o;
  wire [31:0] n9927_data; // mem_rd
  wire [31:0] n9928_data; // mem_rd
  assign addr_out = n1074_o;
  assign data_write = n278_o;
  assign nwr = n78_o;
  assign nuds = n89_o;
  assign nlds = n90_o;
  assign busstate = state;
  assign longword = n56_o;
  assign nresetout = n82_o;
  assign fc = n9925_o;
  assign clr_berr = n98_o;
  assign skipfetch = n9109_o;
  assign regin_out = regin;
  assign cacr_out = cacr;
  assign vbr_out = vbr;
  /* TG68KdotC_Kernel.vhd:148:16  */
  assign use_vbr_stackframe = n9811_q; // (signal)
  /* TG68KdotC_Kernel.vhd:150:16  */
  assign syncreset = n9813_q; // (signal)
  /* TG68KdotC_Kernel.vhd:151:16  */
  assign reset = n9815_q; // (signal)
  /* TG68KdotC_Kernel.vhd:152:16  */
  assign clkena_lw = n94_o; // (signal)
  /* TG68KdotC_Kernel.vhd:153:16  */
  assign tg68_pc = n9816_q; // (signal)
  /* TG68KdotC_Kernel.vhd:154:16  */
  assign tmp_tg68_pc = n9818_q; // (signal)
  /* TG68KdotC_Kernel.vhd:155:16  */
  assign tg68_pc_add = n1175_o; // (signal)
  /* TG68KdotC_Kernel.vhd:156:16  */
  assign pc_dataa = n1081_o; // (signal)
  /* TG68KdotC_Kernel.vhd:157:16  */
  assign pc_datab = n1174_o; // (signal)
  /* TG68KdotC_Kernel.vhd:158:16  */
  assign memaddr = n9820_q; // (signal)
  /* TG68KdotC_Kernel.vhd:159:16  */
  assign state = n9821_q; // (signal)
  /* TG68KdotC_Kernel.vhd:160:16  */
  assign datatype = n9126_o; // (signal)
  /* TG68KdotC_Kernel.vhd:161:16  */
  assign set_datatype = n9127_o; // (signal)
  /* TG68KdotC_Kernel.vhd:162:16  */
  assign exe_datatype = n9822_q; // (signal)
  /* TG68KdotC_Kernel.vhd:163:16  */
  assign setstate = n9169_o; // (signal)
  /* TG68KdotC_Kernel.vhd:164:16  */
  assign setaddrvalue = n9172_o; // (signal)
  /* TG68KdotC_Kernel.vhd:165:16  */
  assign addrvalue = n9823_q; // (signal)
  /* TG68KdotC_Kernel.vhd:167:16  */
  assign opcode = n9824_q; // (signal)
  /* TG68KdotC_Kernel.vhd:168:16  */
  assign exe_opcode = n9825_q; // (signal)
  /* TG68KdotC_Kernel.vhd:169:16  */
  assign sndopc = n9827_q; // (signal)
  /* TG68KdotC_Kernel.vhd:171:16  */
  assign exe_pc = n9828_q; // (signal)
  /* TG68KdotC_Kernel.vhd:172:16  */
  assign last_opc_pc = n9829_q; // (signal)
  /* TG68KdotC_Kernel.vhd:173:16  */
  assign last_opc_read = n9830_q; // (signal)
  /* TG68KdotC_Kernel.vhd:175:16  */
  assign reg_qa = n9928_data; // (signal)
  /* TG68KdotC_Kernel.vhd:176:16  */
  assign reg_qb = n9927_data; // (signal)
  /* TG68KdotC_Kernel.vhd:177:16  */
  assign wwrena = n392_o; // (signal)
  /* TG68KdotC_Kernel.vhd:177:23  */
  assign lwrena = n395_o; // (signal)
  /* TG68KdotC_Kernel.vhd:178:16  */
  assign bwrena = n398_o; // (signal)
  /* TG68KdotC_Kernel.vhd:179:16  */
  assign regwrena_now = n9175_o; // (signal)
  /* TG68KdotC_Kernel.vhd:180:16  */
  assign rf_dest_addr = n440_o; // (signal)
  /* TG68KdotC_Kernel.vhd:181:16  */
  assign rf_source_addr = n478_o; // (signal)
  /* TG68KdotC_Kernel.vhd:182:16  */
  assign rf_source_addrd = n9833_q; // (signal)
  /* TG68KdotC_Kernel.vhd:184:16  */
  assign regin = n9834_o; // (signal)
  /* TG68KdotC_Kernel.vhd:187:16  */
  assign rdindex_a = n9838_q; // (signal)
  /* TG68KdotC_Kernel.vhd:188:16  */
  assign rdindex_b = n9840_q; // (signal)
  /* TG68KdotC_Kernel.vhd:189:16  */
  assign wr_areg = n9842_q; // (signal)
  /* TG68KdotC_Kernel.vhd:192:16  */
  assign addr = n1073_o; // (signal)
  /* TG68KdotC_Kernel.vhd:193:16  */
  assign memaddr_reg = n1077_o; // (signal)
  /* TG68KdotC_Kernel.vhd:194:16  */
  assign memaddr_delta = n1072_o; // (signal)
  /* TG68KdotC_Kernel.vhd:195:16  */
  assign memaddr_delta_rega = n9844_q; // (signal)
  /* TG68KdotC_Kernel.vhd:196:16  */
  assign memaddr_delta_regb = n9846_q; // (signal)
  /* TG68KdotC_Kernel.vhd:197:16  */
  assign use_base = n9848_q; // (signal)
  /* TG68KdotC_Kernel.vhd:199:16  */
  assign ea_data = n9849_q; // (signal)
  /* TG68KdotC_Kernel.vhd:200:16  */
  assign op1out = n494_o; // (signal)
  /* TG68KdotC_Kernel.vhd:201:16  */
  assign op2out = n9850_o; // (signal)
  /* TG68KdotC_Kernel.vhd:202:16  */
  assign op1outbrief = n839_o; // (signal)
  /* TG68KdotC_Kernel.vhd:204:16  */
  assign aluout = alu_n42; // (signal)
  /* TG68KdotC_Kernel.vhd:205:16  */
  assign data_write_tmp = n9852_q; // (signal)
  /* TG68KdotC_Kernel.vhd:206:16  */
  assign data_write_muxin = n241_o; // (signal)
  /* TG68KdotC_Kernel.vhd:207:16  */
  assign data_write_mux = n250_o; // (signal)
  /* TG68KdotC_Kernel.vhd:208:16  */
  assign nextpass = n9853_q; // (signal)
  /* TG68KdotC_Kernel.vhd:209:16  */
  assign setnextpass = n9180_o; // (signal)
  /* TG68KdotC_Kernel.vhd:210:16  */
  assign setdispbyte = n9182_o; // (signal)
  /* TG68KdotC_Kernel.vhd:211:16  */
  assign setdisp = n9192_o; // (signal)
  /* TG68KdotC_Kernel.vhd:212:16  */
  assign regdirectsource = n7810_o; // (signal)
  /* TG68KdotC_Kernel.vhd:213:16  */
  assign addsub_q = alu_n41; // (signal)
  /* TG68KdotC_Kernel.vhd:214:16  */
  assign briefdata = n875_o; // (signal)
  /* TG68KdotC_Kernel.vhd:215:16  */
  assign c_out = alu_n40; // (signal)
  /* TG68KdotC_Kernel.vhd:218:16  */
  assign memaddr_a = n9855_o; // (signal)
  /* TG68KdotC_Kernel.vhd:220:16  */
  assign tg68_pc_brw = n9196_o; // (signal)
  /* TG68KdotC_Kernel.vhd:221:16  */
  assign tg68_pc_word = n9856_q; // (signal)
  /* TG68KdotC_Kernel.vhd:222:16  */
  assign getbrief = n7812_o; // (signal)
  /* TG68KdotC_Kernel.vhd:223:16  */
  assign brief = n9857_q; // (signal)
  /* TG68KdotC_Kernel.vhd:224:16  */
  assign data_is_source = n7814_o; // (signal)
  /* TG68KdotC_Kernel.vhd:225:16  */
  assign store_in_tmp = n9858_q; // (signal)
  /* TG68KdotC_Kernel.vhd:226:16  */
  assign write_back = n8096_o; // (signal)
  /* TG68KdotC_Kernel.vhd:227:16  */
  assign exec_write_back = n9859_q; // (signal)
  /* TG68KdotC_Kernel.vhd:228:16  */
  assign setstackaddr = n9214_o; // (signal)
  /* TG68KdotC_Kernel.vhd:229:16  */
  assign writepc = n9216_o; // (signal)
  /* TG68KdotC_Kernel.vhd:230:16  */
  assign writepcbig = n9860_q; // (signal)
  /* TG68KdotC_Kernel.vhd:231:16  */
  assign set_writepcbig = n9219_o; // (signal)
  /* TG68KdotC_Kernel.vhd:232:16  */
  assign writepcnext = n9861_q; // (signal)
  /* TG68KdotC_Kernel.vhd:233:16  */
  assign setopcode = n1211_o; // (signal)
  /* TG68KdotC_Kernel.vhd:234:16  */
  assign decodeopc = n9862_q; // (signal)
  /* TG68KdotC_Kernel.vhd:235:16  */
  assign execopc = n9863_q; // (signal)
  /* TG68KdotC_Kernel.vhd:236:16  */
  assign execopc_alu = n60_o; // (signal)
  /* TG68KdotC_Kernel.vhd:237:16  */
  assign setexecopc = n1236_o; // (signal)
  /* TG68KdotC_Kernel.vhd:238:16  */
  assign endopc = n9864_q; // (signal)
  /* TG68KdotC_Kernel.vhd:239:16  */
  assign setendopc = n1215_o; // (signal)
  /* TG68KdotC_Kernel.vhd:240:16  */
  assign flags = alu_n39; // (signal)
  /* TG68KdotC_Kernel.vhd:241:16  */
  assign flagssr = n9865_q; // (signal)
  /* TG68KdotC_Kernel.vhd:242:16  */
  assign srin = n1785_o; // (signal)
  /* TG68KdotC_Kernel.vhd:243:16  */
  assign exec_direct = n9866_q; // (signal)
  /* TG68KdotC_Kernel.vhd:244:16  */
  assign exec_tas = n9868_q; // (signal)
  /* TG68KdotC_Kernel.vhd:245:16  */
  assign set_exec_tas = n7824_o; // (signal)
  /* TG68KdotC_Kernel.vhd:247:16  */
  assign exe_condition = n9643_o; // (signal)
  /* TG68KdotC_Kernel.vhd:248:16  */
  assign ea_only = n7827_o; // (signal)
  /* TG68KdotC_Kernel.vhd:249:16  */
  assign source_areg = n9222_o; // (signal)
  /* TG68KdotC_Kernel.vhd:250:16  */
  assign source_lowbits = n8098_o; // (signal)
  /* TG68KdotC_Kernel.vhd:251:16  */
  assign source_ldrlbits = n9225_o; // (signal)
  /* TG68KdotC_Kernel.vhd:252:16  */
  assign source_ldrmbits = n9229_o; // (signal)
  /* TG68KdotC_Kernel.vhd:253:16  */
  assign source_2ndhbits = n7836_o; // (signal)
  /* TG68KdotC_Kernel.vhd:254:16  */
  assign source_2ndmbits = n9233_o; // (signal)
  /* TG68KdotC_Kernel.vhd:255:16  */
  assign source_2ndlbits = n9236_o; // (signal)
  /* TG68KdotC_Kernel.vhd:256:16  */
  assign dest_areg = n9241_o; // (signal)
  /* TG68KdotC_Kernel.vhd:257:16  */
  assign dest_ldrareg = n9243_o; // (signal)
  /* TG68KdotC_Kernel.vhd:258:16  */
  assign dest_ldrhbits = n9248_o; // (signal)
  /* TG68KdotC_Kernel.vhd:259:16  */
  assign dest_ldrlbits = n9251_o; // (signal)
  /* TG68KdotC_Kernel.vhd:260:16  */
  assign dest_2ndhbits = n9257_o; // (signal)
  /* TG68KdotC_Kernel.vhd:261:16  */
  assign dest_2ndlbits = n9261_o; // (signal)
  /* TG68KdotC_Kernel.vhd:262:16  */
  assign dest_hbits = n9266_o; // (signal)
  /* TG68KdotC_Kernel.vhd:263:16  */
  assign rot_bits = n9869_q; // (signal)
  /* TG68KdotC_Kernel.vhd:264:16  */
  assign set_rot_bits = n7850_o; // (signal)
  /* TG68KdotC_Kernel.vhd:265:16  */
  assign rot_cnt = n9870_q; // (signal)
  /* TG68KdotC_Kernel.vhd:266:16  */
  assign set_rot_cnt = n9267_o; // (signal)
  /* TG68KdotC_Kernel.vhd:267:16  */
  assign movem_actiond = n9872_q; // (signal)
  /* TG68KdotC_Kernel.vhd:268:16  */
  assign movem_regaddr = n9873_o; // (signal)
  /* TG68KdotC_Kernel.vhd:269:16  */
  assign movem_mux = n9785_o; // (signal)
  /* TG68KdotC_Kernel.vhd:270:16  */
  assign movem_presub = n7853_o; // (signal)
  /* TG68KdotC_Kernel.vhd:271:16  */
  assign movem_run = n9787_o; // (signal)
  /* TG68KdotC_Kernel.vhd:273:16  */
  assign set_direct_data = n9271_o; // (signal)
  /* TG68KdotC_Kernel.vhd:274:16  */
  assign use_direct_data = n9875_q; // (signal)
  /* TG68KdotC_Kernel.vhd:275:16  */
  assign direct_data = n9876_q; // (signal)
  /* TG68KdotC_Kernel.vhd:277:16  */
  assign set_v_flag = alu_n38; // (signal)
  /* TG68KdotC_Kernel.vhd:278:16  */
  assign set_vectoraddr = n9274_o; // (signal)
  /* TG68KdotC_Kernel.vhd:279:16  */
  assign writesr = n9278_o; // (signal)
  /* TG68KdotC_Kernel.vhd:280:16  */
  assign trap_berr = n9877_q; // (signal)
  /* TG68KdotC_Kernel.vhd:281:16  */
  assign trap_illegal = n9280_o; // (signal)
  /* TG68KdotC_Kernel.vhd:282:16  */
  assign trap_addr_error = n7861_o; // (signal)
  /* TG68KdotC_Kernel.vhd:283:16  */
  assign trap_priv = n7864_o; // (signal)
  /* TG68KdotC_Kernel.vhd:284:16  */
  assign trap_trace = n9878_q; // (signal)
  /* TG68KdotC_Kernel.vhd:285:16  */
  assign trap_1010 = n7867_o; // (signal)
  /* TG68KdotC_Kernel.vhd:286:16  */
  assign trap_1111 = n7870_o; // (signal)
  /* TG68KdotC_Kernel.vhd:287:16  */
  assign trap_trap = n7873_o; // (signal)
  /* TG68KdotC_Kernel.vhd:288:16  */
  assign trap_trapv = n7876_o; // (signal)
  /* TG68KdotC_Kernel.vhd:289:16  */
  assign trap_interrupt = n9879_q; // (signal)
  /* TG68KdotC_Kernel.vhd:290:16  */
  assign trapmake = n9281_o; // (signal)
  /* TG68KdotC_Kernel.vhd:291:16  */
  assign trapd = n9880_q; // (signal)
  /* TG68KdotC_Kernel.vhd:292:16  */
  assign trap_sr = n9881_q; // (signal)
  /* TG68KdotC_Kernel.vhd:293:16  */
  assign make_trace = n9882_q; // (signal)
  /* TG68KdotC_Kernel.vhd:294:16  */
  assign make_berr = n9883_q; // (signal)
  /* TG68KdotC_Kernel.vhd:295:16  */
  assign usestackframe2 = n9884_q; // (signal)
  /* TG68KdotC_Kernel.vhd:297:16  */
  assign set_stop = n7882_o; // (signal)
  /* TG68KdotC_Kernel.vhd:298:16  */
  assign stop = n9885_q; // (signal)
  /* TG68KdotC_Kernel.vhd:299:16  */
  assign trap_vector = n9887_q; // (signal)
  /* TG68KdotC_Kernel.vhd:300:16  */
  assign trap_vector_vbr = n917_o; // (signal)
  /* TG68KdotC_Kernel.vhd:301:16  */
  assign usp = n9889_q; // (signal)
  /* TG68KdotC_Kernel.vhd:306:16  */
  assign ipl_nr = n1238_o; // (signal)
  /* TG68KdotC_Kernel.vhd:307:16  */
  assign ripl_nr = n9890_q; // (signal)
  /* TG68KdotC_Kernel.vhd:308:16  */
  assign ipl_vec = n9891_q; // (signal)
  /* TG68KdotC_Kernel.vhd:309:16  */
  assign interrupt = n9892_q; // (signal)
  /* TG68KdotC_Kernel.vhd:310:16  */
  assign setinterrupt = n1218_o; // (signal)
  /* TG68KdotC_Kernel.vhd:311:16  */
  assign svmode = n9893_q; // (signal)
  /* TG68KdotC_Kernel.vhd:312:16  */
  assign presvmode = n9894_q; // (signal)
  /* TG68KdotC_Kernel.vhd:313:16  */
  assign suppress_base = n9895_q; // (signal)
  /* TG68KdotC_Kernel.vhd:314:16  */
  assign set_suppress_base = n9284_o; // (signal)
  /* TG68KdotC_Kernel.vhd:315:16  */
  assign set_z_error = n9286_o; // (signal)
  /* TG68KdotC_Kernel.vhd:316:16  */
  assign z_error = n9896_q; // (signal)
  /* TG68KdotC_Kernel.vhd:317:16  */
  assign ea_build_now = n8035_o; // (signal)
  /* TG68KdotC_Kernel.vhd:318:16  */
  assign build_logical = n7888_o; // (signal)
  /* TG68KdotC_Kernel.vhd:319:16  */
  assign build_bcd = n7891_o; // (signal)
  /* TG68KdotC_Kernel.vhd:321:16  */
  assign data_read = n9897_o; // (signal)
  /* TG68KdotC_Kernel.vhd:322:16  */
  assign bf_ext_in = n9899_q; // (signal)
  /* TG68KdotC_Kernel.vhd:323:16  */
  assign bf_ext_out = alu_n36; // (signal)
  /* TG68KdotC_Kernel.vhd:325:16  */
  assign long_start = n234_o; // (signal)
  /* TG68KdotC_Kernel.vhd:326:16  */
  assign long_start_alu = n58_o; // (signal)
  /* TG68KdotC_Kernel.vhd:327:16  */
  assign non_aligned = n72_o; // (signal)
  /* TG68KdotC_Kernel.vhd:328:16  */
  assign check_aligned = n7894_o; // (signal)
  /* TG68KdotC_Kernel.vhd:329:16  */
  assign long_done = n236_o; // (signal)
  /* TG68KdotC_Kernel.vhd:330:16  */
  assign memmask = n9900_q; // (signal)
  /* TG68KdotC_Kernel.vhd:331:16  */
  assign set_memmask = n1769_o; // (signal)
  /* TG68KdotC_Kernel.vhd:332:16  */
  assign memread = n9901_q; // (signal)
  /* TG68KdotC_Kernel.vhd:333:16  */
  assign wbmemmask = n9902_q; // (signal)
  /* TG68KdotC_Kernel.vhd:334:16  */
  assign memmaskmux = n85_o; // (signal)
  /* TG68KdotC_Kernel.vhd:335:16  */
  assign oddout = n9903_q; // (signal)
  /* TG68KdotC_Kernel.vhd:336:16  */
  assign set_oddout = n1694_o; // (signal)
  /* TG68KdotC_Kernel.vhd:337:16  */
  assign pcbase = n9904_q; // (signal)
  /* TG68KdotC_Kernel.vhd:338:16  */
  assign set_pcbase = n2160_o; // (signal)
  /* TG68KdotC_Kernel.vhd:340:16  */
  assign last_data_read = n9905_q; // (signal)
  /* TG68KdotC_Kernel.vhd:341:16  */
  assign last_data_in = n9906_q; // (signal)
  /* TG68KdotC_Kernel.vhd:343:16  */
  assign bf_offset = n9907_o; // (signal)
  /* TG68KdotC_Kernel.vhd:344:16  */
  assign bf_width = n9908_o; // (signal)
  /* TG68KdotC_Kernel.vhd:345:16  */
  assign bf_bhits = n1692_o; // (signal)
  /* TG68KdotC_Kernel.vhd:346:16  */
  assign bf_shift = n1749_o; // (signal)
  /* TG68KdotC_Kernel.vhd:347:16  */
  assign alu_width = n9909_q; // (signal)
  /* TG68KdotC_Kernel.vhd:348:16  */
  assign alu_bf_shift = n9910_q; // (signal)
  /* TG68KdotC_Kernel.vhd:349:16  */
  assign bf_loffset = n9911_o; // (signal)
  /* TG68KdotC_Kernel.vhd:350:16  */
  assign bf_full_offset = n1682_o; // (signal)
  /* TG68KdotC_Kernel.vhd:351:16  */
  assign alu_bf_ffo_offset = n9912_q; // (signal)
  /* TG68KdotC_Kernel.vhd:352:16  */
  assign alu_bf_loffset = n9913_q; // (signal)
  /* TG68KdotC_Kernel.vhd:354:16  */
  assign movec_data = n9538_o; // (signal)
  /* TG68KdotC_Kernel.vhd:355:16  */
  assign vbr = n9914_q; // (signal)
  /* TG68KdotC_Kernel.vhd:356:16  */
  assign cacr = n9915_q; // (signal)
  /* TG68KdotC_Kernel.vhd:357:16  */
  assign dfc = n9916_q; // (signal)
  /* TG68KdotC_Kernel.vhd:358:16  */
  assign sfc = n9917_q; // (signal)
  /* TG68KdotC_Kernel.vhd:361:16  */
  assign set = n9918_o; // (signal)
  /* TG68KdotC_Kernel.vhd:362:16  */
  assign set_exec = n9919_o; // (signal)
  /* TG68KdotC_Kernel.vhd:363:16  */
  assign exec = n9921_q; // (signal)
  /* TG68KdotC_Kernel.vhd:365:16  */
  assign micro_state = n9922_q; // (signal)
  /* TG68KdotC_Kernel.vhd:366:16  */
  assign next_micro_state = n9473_o; // (signal)
  /* TG68KdotC_Kernel.vhd:405:49  */
  assign n34_o = last_data_read[15:0];
  /* TG68KdotC_Kernel.vhd:406:39  */
  assign n35_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:410:31  */
  assign alu_n36 = alu_bf_ext_out; // (signal)
  /* TG68KdotC_Kernel.vhd:414:45  */
  assign n37_o = alu_bf_loffset[4:0];
  /* TG68KdotC_Kernel.vhd:416:31  */
  assign alu_n38 = alu_set_v_flag; // (signal)
  /* TG68KdotC_Kernel.vhd:417:26  */
  assign alu_n39 = alu_flags; // (signal)
  /* TG68KdotC_Kernel.vhd:418:26  */
  assign alu_n40 = alu_c_out; // (signal)
  /* TG68KdotC_Kernel.vhd:419:29  */
  assign alu_n41 = alu_addsub_q; // (signal)
  /* TG68KdotC_Kernel.vhd:420:27  */
  assign alu_n42 = alu_aluout; // (signal)
  /* TG68KdotC_Kernel.vhd:372:1  */
  tg68k_alu_2_1_2_1 alu (
    .clk(clk),
    .reset(reset),
    .clkena_lw(clkena_lw),
    .cpu(cpu),
    .execopc(execopc_alu),
    .decodeopc(decodeopc),
    .exe_condition(exe_condition),
    .exec_tas(exec_tas),
    .long_start(long_start_alu),
    .non_aligned(non_aligned),
    .check_aligned(check_aligned),
    .movem_presub(movem_presub),
    .set_stop(set_stop),
    .z_error(z_error),
    .rot_bits(rot_bits),
    .exec(exec),
    .op1out(op1out),
    .op2out(op2out),
    .reg_qa(reg_qa),
    .reg_qb(reg_qb),
    .opcode(opcode),
    .exe_opcode(exe_opcode),
    .exe_datatype(exe_datatype),
    .sndopc(sndopc),
    .last_data_read(n34_o),
    .data_read(n35_o),
    .flagssr(flagssr),
    .micro_state(micro_state),
    .bf_ext_in(bf_ext_in),
    .bf_shift(alu_bf_shift),
    .bf_width(alu_width),
    .bf_ffo_offset(alu_bf_ffo_offset),
    .bf_loffset(n37_o),
    .bf_ext_out(alu_bf_ext_out),
    .set_v_flag(alu_set_v_flag),
    .flags(alu_flags),
    .c_out(alu_c_out),
    .addsub_q(alu_addsub_q),
    .aluout(alu_aluout));
  /* TG68KdotC_Kernel.vhd:424:35  */
  assign n55_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:424:21  */
  assign n56_o = ~n55_o;
  /* TG68KdotC_Kernel.vhd:426:48  */
  assign n57_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:426:34  */
  assign n58_o = ~n57_o;
  /* TG68KdotC_Kernel.vhd:427:39  */
  assign n59_o = exec[84];
  /* TG68KdotC_Kernel.vhd:427:32  */
  assign n60_o = execopc | n59_o;
  /* TG68KdotC_Kernel.vhd:431:31  */
  assign n63_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:431:44  */
  assign n65_o = n63_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:431:66  */
  assign n66_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:431:79  */
  assign n68_o = n66_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:431:52  */
  assign n69_o = n65_o | n68_o;
  /* TG68KdotC_Kernel.vhd:431:17  */
  assign n72_o = n69_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:441:30  */
  assign n77_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:441:20  */
  assign n78_o = n77_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:443:35  */
  assign n81_o = exec[74];
  /* TG68KdotC_Kernel.vhd:443:26  */
  assign n82_o = n81_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:447:40  */
  assign n84_o = addr[0];
  /* TG68KdotC_Kernel.vhd:447:31  */
  assign n85_o = n84_o ? memmask : n88_o;
  /* TG68KdotC_Kernel.vhd:447:62  */
  assign n86_o = memmask[4:0];
  /* TG68KdotC_Kernel.vhd:447:75  */
  assign n88_o = {n86_o, 1'b1};
  /* TG68KdotC_Kernel.vhd:448:27  */
  assign n89_o = memmaskmux[5];
  /* TG68KdotC_Kernel.vhd:449:27  */
  assign n90_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:450:59  */
  assign n92_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:450:45  */
  assign n93_o = n92_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:450:26  */
  assign n94_o = n93_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:451:44  */
  assign n97_o = trap_berr & setopcode;
  /* TG68KdotC_Kernel.vhd:451:25  */
  assign n98_o = n97_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:455:26  */
  assign n102_o = ~nreset;
  /* TG68KdotC_Kernel.vhd:460:55  */
  assign n104_o = syncreset[2:0];
  /* TG68KdotC_Kernel.vhd:460:67  */
  assign n106_o = {n104_o, 1'b1};
  /* TG68KdotC_Kernel.vhd:461:55  */
  assign n107_o = syncreset[3];
  /* TG68KdotC_Kernel.vhd:461:42  */
  assign n108_o = ~n107_o;
  /* TG68KdotC_Kernel.vhd:465:52  */
  assign n118_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:465:60  */
  assign n120_o = 1'b1 & n118_o;
  /* TG68KdotC_Kernel.vhd:465:45  */
  assign n122_o = 1'b0 | n120_o;
  /* TG68KdotC_Kernel.vhd:465:25  */
  assign n125_o = n122_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:475:30  */
  assign n130_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:475:33  */
  assign n131_o = ~n130_o;
  /* TG68KdotC_Kernel.vhd:476:50  */
  assign n132_o = last_data_in[15:0];
  /* TG68KdotC_Kernel.vhd:476:63  */
  assign n133_o = {n132_o, data_in};
  /* TG68KdotC_Kernel.vhd:478:50  */
  assign n134_o = last_data_in[23:0];
  /* TG68KdotC_Kernel.vhd:478:71  */
  assign n135_o = data_in[15:8];
  /* TG68KdotC_Kernel.vhd:478:63  */
  assign n136_o = {n134_o, n135_o};
  /* TG68KdotC_Kernel.vhd:480:27  */
  assign n138_o = memread[0];
  /* TG68KdotC_Kernel.vhd:480:46  */
  assign n139_o = memread[1:0];
  /* TG68KdotC_Kernel.vhd:480:58  */
  assign n141_o = n139_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:480:78  */
  assign n142_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:480:64  */
  assign n143_o = n142_o & n141_o;
  /* TG68KdotC_Kernel.vhd:480:35  */
  assign n144_o = n138_o | n143_o;
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n145_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n146_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n147_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n148_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n149_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n150_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n151_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n152_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n153_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n154_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n155_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n156_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n157_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n158_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n159_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n160_o = data_read[15];
  assign n161_o = {n145_o, n146_o, n147_o, n148_o};
  assign n162_o = {n149_o, n150_o, n151_o, n152_o};
  assign n163_o = {n153_o, n154_o, n155_o, n156_o};
  assign n164_o = {n157_o, n158_o, n159_o, n160_o};
  assign n165_o = {n161_o, n162_o, n163_o, n164_o};
  assign n166_o = n133_o[31:16];
  assign n167_o = n136_o[31:16];
  /* TG68KdotC_Kernel.vhd:475:17  */
  assign n168_o = n131_o ? n166_o : n167_o;
  /* TG68KdotC_Kernel.vhd:480:17  */
  assign n169_o = n144_o ? n165_o : n168_o;
  assign n170_o = n133_o[15:0];
  assign n171_o = n136_o[15:0];
  /* TG68KdotC_Kernel.vhd:475:17  */
  assign n172_o = n131_o ? n170_o : n171_o;
  /* TG68KdotC_Kernel.vhd:485:51  */
  assign n175_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:485:42  */
  assign n176_o = n175_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:486:46  */
  assign n177_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:486:49  */
  assign n178_o = ~n177_o;
  /* TG68KdotC_Kernel.vhd:487:66  */
  assign n179_o = last_data_in[23:16];
  /* TG68KdotC_Kernel.vhd:489:66  */
  assign n180_o = last_data_in[31:24];
  /* TG68KdotC_Kernel.vhd:486:33  */
  assign n181_o = n178_o ? n179_o : n180_o;
  /* TG68KdotC_Kernel.vhd:495:41  */
  assign n184_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:495:54  */
  assign n185_o = exec[38];
  /* TG68KdotC_Kernel.vhd:495:47  */
  assign n186_o = n184_o | n185_o;
  /* TG68KdotC_Kernel.vhd:497:49  */
  assign n187_o = state[1];
  /* TG68KdotC_Kernel.vhd:497:52  */
  assign n188_o = ~n187_o;
  /* TG68KdotC_Kernel.vhd:497:68  */
  assign n189_o = memmask[1];
  /* TG68KdotC_Kernel.vhd:497:71  */
  assign n190_o = ~n189_o;
  /* TG68KdotC_Kernel.vhd:497:57  */
  assign n191_o = n190_o & n188_o;
  /* TG68KdotC_Kernel.vhd:499:52  */
  assign n192_o = state[1];
  /* TG68KdotC_Kernel.vhd:499:55  */
  assign n193_o = ~n192_o;
  /* TG68KdotC_Kernel.vhd:499:70  */
  assign n194_o = memread[1];
  /* TG68KdotC_Kernel.vhd:499:60  */
  assign n195_o = n193_o | n194_o;
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n196_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n197_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n198_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n199_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n200_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n201_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n202_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n203_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n204_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n205_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n206_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n207_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n208_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n209_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n210_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n211_o = data_in[15];
  assign n212_o = {n196_o, n197_o, n198_o, n199_o};
  assign n213_o = {n200_o, n201_o, n202_o, n203_o};
  assign n214_o = {n204_o, n205_o, n206_o, n207_o};
  assign n215_o = {n208_o, n209_o, n210_o, n211_o};
  assign n216_o = {n212_o, n213_o, n214_o, n215_o};
  assign n217_o = data_read[31:16];
  /* TG68KdotC_Kernel.vhd:499:41  */
  assign n218_o = n195_o ? n216_o : n217_o;
  /* TG68KdotC_Kernel.vhd:497:41  */
  assign n219_o = n191_o ? last_opc_read : n218_o;
  assign n220_o = data_read[15:0];
  assign n221_o = {n219_o, n220_o};
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n222_o = n225_o ? n221_o : last_data_read;
  /* TG68KdotC_Kernel.vhd:503:61  */
  assign n223_o = last_data_in[15:0];
  /* TG68KdotC_Kernel.vhd:503:74  */
  assign n224_o = {n223_o, data_in};
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n225_o = n186_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n226_o = clkena_in ? n224_o : last_data_in;
  /* TG68KdotC_Kernel.vhd:492:25  */
  assign n228_o = reset ? 32'b00000000000000000000000000000000 : n222_o;
  /* TG68KdotC_Kernel.vhd:492:25  */
  assign n229_o = reset ? last_data_in : n226_o;
  /* TG68KdotC_Kernel.vhd:507:65  */
  assign n233_o = memmask[1];
  /* TG68KdotC_Kernel.vhd:507:54  */
  assign n234_o = ~n233_o;
  /* TG68KdotC_Kernel.vhd:508:64  */
  assign n235_o = memread[1];
  /* TG68KdotC_Kernel.vhd:508:53  */
  assign n236_o = ~n235_o;
  /* TG68KdotC_Kernel.vhd:514:24  */
  assign n240_o = exec[40];
  /* TG68KdotC_Kernel.vhd:514:17  */
  assign n241_o = n240_o ? reg_qb : data_write_tmp;
  /* TG68KdotC_Kernel.vhd:527:39  */
  assign n242_o = addr[0];
  /* TG68KdotC_Kernel.vhd:527:34  */
  assign n243_o = oddout == n242_o;
  /* TG68KdotC_Kernel.vhd:528:61  */
  assign n245_o = {8'bX, bf_ext_out};
  /* TG68KdotC_Kernel.vhd:528:72  */
  assign n246_o = {n245_o, data_write_muxin};
  /* TG68KdotC_Kernel.vhd:530:61  */
  assign n247_o = {bf_ext_out, data_write_muxin};
  /* TG68KdotC_Kernel.vhd:530:78  */
  assign n249_o = {n247_o, 8'bX};
  /* TG68KdotC_Kernel.vhd:527:25  */
  assign n250_o = n243_o ? n246_o : n249_o;
  /* TG68KdotC_Kernel.vhd:534:30  */
  assign n251_o = memmaskmux[1];
  /* TG68KdotC_Kernel.vhd:534:33  */
  assign n252_o = ~n251_o;
  /* TG68KdotC_Kernel.vhd:535:53  */
  assign n253_o = data_write_mux[47:32];
  /* TG68KdotC_Kernel.vhd:536:33  */
  assign n254_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:536:36  */
  assign n255_o = ~n254_o;
  /* TG68KdotC_Kernel.vhd:537:53  */
  assign n256_o = data_write_mux[31:16];
  /* TG68KdotC_Kernel.vhd:540:38  */
  assign n257_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:540:51  */
  assign n259_o = n257_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:541:61  */
  assign n260_o = data_write_mux[7:0];
  /* TG68KdotC_Kernel.vhd:541:90  */
  assign n261_o = data_write_mux[7:0];
  /* TG68KdotC_Kernel.vhd:541:74  */
  assign n262_o = {n260_o, n261_o};
  /* TG68KdotC_Kernel.vhd:542:41  */
  assign n263_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:542:54  */
  assign n265_o = n263_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:543:61  */
  assign n266_o = data_write_mux[15:8];
  /* TG68KdotC_Kernel.vhd:543:91  */
  assign n267_o = data_write_mux[15:8];
  /* TG68KdotC_Kernel.vhd:543:75  */
  assign n268_o = {n266_o, n267_o};
  /* TG68KdotC_Kernel.vhd:545:61  */
  assign n269_o = data_write_mux[15:0];
  /* TG68KdotC_Kernel.vhd:542:25  */
  assign n270_o = n265_o ? n268_o : n269_o;
  /* TG68KdotC_Kernel.vhd:540:25  */
  assign n271_o = n259_o ? n262_o : n270_o;
  /* TG68KdotC_Kernel.vhd:536:17  */
  assign n272_o = n255_o ? n256_o : n271_o;
  /* TG68KdotC_Kernel.vhd:534:17  */
  assign n273_o = n252_o ? n253_o : n272_o;
  /* TG68KdotC_Kernel.vhd:548:24  */
  assign n274_o = exec[72];
  /* TG68KdotC_Kernel.vhd:549:53  */
  assign n275_o = data_write_tmp[15:8];
  /* TG68KdotC_Kernel.vhd:549:83  */
  assign n276_o = data_write_tmp[15:8];
  /* TG68KdotC_Kernel.vhd:549:67  */
  assign n277_o = {n275_o, n276_o};
  /* TG68KdotC_Kernel.vhd:548:17  */
  assign n278_o = n274_o ? n277_o : n273_o;
  /* TG68KdotC_Kernel.vhd:563:56  */
  assign n291_o = rf_dest_addr[3];
  /* TG68KdotC_Kernel.vhd:570:40  */
  assign n299_o = exec[65];
  /* TG68KdotC_Kernel.vhd:561:21  */
  assign n302_o = wwrena & clkena_lw;
  /* TG68KdotC_Kernel.vhd:561:21  */
  assign n306_o = n299_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:583:24  */
  assign n316_o = exec[30];
  /* TG68KdotC_Kernel.vhd:585:27  */
  assign n317_o = exec[62];
  /* TG68KdotC_Kernel.vhd:585:44  */
  assign n318_o = ea_only & n317_o;
  /* TG68KdotC_Kernel.vhd:587:27  */
  assign n319_o = exec[66];
  /* TG68KdotC_Kernel.vhd:589:27  */
  assign n320_o = exec[32];
  /* TG68KdotC_Kernel.vhd:594:53  */
  assign n325_o = reg_qa[15:8];
  assign n326_o = memaddr[15:8];
  assign n327_o = memaddr_a[15:8];
  assign n328_o = usp[15:8];
  assign n329_o = movec_data[15:8];
  assign n330_o = aluout[15:8];
  /* TG68KdotC_Kernel.vhd:589:17  */
  assign n331_o = n320_o ? n329_o : n330_o;
  /* TG68KdotC_Kernel.vhd:587:17  */
  assign n332_o = n319_o ? n328_o : n331_o;
  /* TG68KdotC_Kernel.vhd:585:17  */
  assign n333_o = n318_o ? n327_o : n332_o;
  /* TG68KdotC_Kernel.vhd:583:17  */
  assign n334_o = n316_o ? n326_o : n333_o;
  /* TG68KdotC_Kernel.vhd:593:17  */
  assign n335_o = bwrena ? n325_o : n334_o;
  assign n336_o = memaddr[31:16];
  assign n337_o = memaddr_a[31:16];
  assign n338_o = usp[31:16];
  assign n339_o = movec_data[31:16];
  assign n340_o = aluout[31:16];
  /* TG68KdotC_Kernel.vhd:589:17  */
  assign n341_o = n320_o ? n339_o : n340_o;
  /* TG68KdotC_Kernel.vhd:587:17  */
  assign n342_o = n319_o ? n338_o : n341_o;
  /* TG68KdotC_Kernel.vhd:585:17  */
  assign n343_o = n318_o ? n337_o : n342_o;
  /* TG68KdotC_Kernel.vhd:583:17  */
  assign n344_o = n316_o ? n336_o : n343_o;
  assign n345_o = memaddr[7:0];
  assign n346_o = memaddr_a[7:0];
  assign n347_o = usp[7:0];
  assign n348_o = movec_data[7:0];
  assign n349_o = aluout[7:0];
  /* TG68KdotC_Kernel.vhd:589:17  */
  assign n350_o = n320_o ? n348_o : n349_o;
  /* TG68KdotC_Kernel.vhd:587:17  */
  assign n351_o = n319_o ? n347_o : n350_o;
  /* TG68KdotC_Kernel.vhd:585:17  */
  assign n352_o = n318_o ? n346_o : n351_o;
  /* TG68KdotC_Kernel.vhd:583:17  */
  assign n353_o = n316_o ? n345_o : n352_o;
  /* TG68KdotC_Kernel.vhd:596:26  */
  assign n354_o = ~lwrena;
  /* TG68KdotC_Kernel.vhd:597:54  */
  assign n355_o = reg_qa[31:16];
  /* TG68KdotC_Kernel.vhd:596:17  */
  assign n356_o = n354_o ? n355_o : n344_o;
  /* TG68KdotC_Kernel.vhd:603:24  */
  assign n357_o = exec[47];
  /* TG68KdotC_Kernel.vhd:603:44  */
  assign n358_o = exec[46];
  /* TG68KdotC_Kernel.vhd:603:37  */
  assign n359_o = n357_o | n358_o;
  /* TG68KdotC_Kernel.vhd:603:65  */
  assign n360_o = exec[41];
  /* TG68KdotC_Kernel.vhd:603:58  */
  assign n361_o = n359_o | n360_o;
  /* TG68KdotC_Kernel.vhd:608:27  */
  assign n362_o = exec[34];
  /* TG68KdotC_Kernel.vhd:611:33  */
  assign n364_o = exe_datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:614:56  */
  assign n365_o = wr_areg | movem_actiond;
  /* TG68KdotC_Kernel.vhd:614:41  */
  assign n368_o = n365_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:613:33  */
  assign n370_o = exe_datatype == 2'b01;
  assign n371_o = {n370_o, n364_o};
  /* TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n371_o)
      2'b10: n374_o = n368_o;
      2'b01: n374_o = 1'b0;
      default: n374_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n371_o)
      2'b10: n377_o = 1'b0;
      2'b01: n377_o = 1'b1;
      default: n377_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n380_o = n362_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n382_o = n362_o ? n374_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n384_o = n362_o ? n377_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n386_o = regwrena_now ? 1'b1 : n380_o;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n388_o = regwrena_now ? 1'b0 : n382_o;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n390_o = regwrena_now ? 1'b0 : n384_o;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n392_o = n361_o ? 1'b1 : n386_o;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n395_o = n361_o ? 1'b1 : n388_o;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n398_o = n361_o ? 1'b0 : n390_o;
  /* TG68KdotC_Kernel.vhd:628:24  */
  assign n403_o = exec[69];
  /* TG68KdotC_Kernel.vhd:630:26  */
  assign n404_o = set[70];
  /* TG68KdotC_Kernel.vhd:631:46  */
  assign n405_o = brief[15:12];
  /* TG68KdotC_Kernel.vhd:632:26  */
  assign n406_o = set[29];
  /* TG68KdotC_Kernel.vhd:634:59  */
  assign n407_o = sndopc[8:6];
  /* TG68KdotC_Kernel.vhd:634:52  */
  assign n409_o = {1'b0, n407_o};
  /* TG68KdotC_Kernel.vhd:639:60  */
  assign n410_o = sndopc[14:12];
  /* TG68KdotC_Kernel.vhd:639:53  */
  assign n411_o = {dest_ldrareg, n410_o};
  /* TG68KdotC_Kernel.vhd:641:55  */
  assign n412_o = last_data_read[15:12];
  /* TG68KdotC_Kernel.vhd:643:59  */
  assign n413_o = last_data_read[2:0];
  /* TG68KdotC_Kernel.vhd:643:44  */
  assign n415_o = {1'b0, n413_o};
  /* TG68KdotC_Kernel.vhd:645:51  */
  assign n416_o = sndopc[2:0];
  /* TG68KdotC_Kernel.vhd:645:44  */
  assign n418_o = {1'b0, n416_o};
  /* TG68KdotC_Kernel.vhd:649:57  */
  assign n419_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:649:50  */
  assign n420_o = {dest_areg, n419_o};
  /* TG68KdotC_Kernel.vhd:651:34  */
  assign n421_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:651:46  */
  assign n423_o = n421_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:651:53  */
  assign n424_o = n423_o | data_is_source;
  /* TG68KdotC_Kernel.vhd:652:65  */
  assign n425_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:652:58  */
  assign n426_o = {dest_areg, n425_o};
  /* TG68KdotC_Kernel.vhd:654:59  */
  assign n427_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:654:52  */
  assign n429_o = {1'b1, n427_o};
  /* TG68KdotC_Kernel.vhd:651:25  */
  assign n430_o = n424_o ? n426_o : n429_o;
  /* TG68KdotC_Kernel.vhd:648:17  */
  assign n431_o = dest_hbits ? n420_o : n430_o;
  /* TG68KdotC_Kernel.vhd:646:17  */
  assign n433_o = setstackaddr ? 4'b1111 : n431_o;
  /* TG68KdotC_Kernel.vhd:644:17  */
  assign n434_o = dest_2ndlbits ? n418_o : n433_o;
  /* TG68KdotC_Kernel.vhd:642:17  */
  assign n435_o = dest_ldrlbits ? n415_o : n434_o;
  /* TG68KdotC_Kernel.vhd:640:17  */
  assign n436_o = dest_ldrhbits ? n412_o : n435_o;
  /* TG68KdotC_Kernel.vhd:638:17  */
  assign n437_o = dest_2ndhbits ? n411_o : n436_o;
  /* TG68KdotC_Kernel.vhd:632:17  */
  assign n438_o = n406_o ? n409_o : n437_o;
  /* TG68KdotC_Kernel.vhd:630:17  */
  assign n439_o = n404_o ? n405_o : n438_o;
  /* TG68KdotC_Kernel.vhd:628:17  */
  assign n440_o = n403_o ? rf_source_addrd : n439_o;
  /* TG68KdotC_Kernel.vhd:664:24  */
  assign n444_o = exec[69];
  /* TG68KdotC_Kernel.vhd:664:49  */
  assign n445_o = set[69];
  /* TG68KdotC_Kernel.vhd:664:43  */
  assign n446_o = n444_o | n445_o;
  /* TG68KdotC_Kernel.vhd:666:65  */
  assign n448_o = movem_regaddr ^ 4'b1111;
  /* TG68KdotC_Kernel.vhd:665:25  */
  assign n449_o = movem_presub ? n448_o : movem_regaddr;
  /* TG68KdotC_Kernel.vhd:671:53  */
  assign n450_o = sndopc[2:0];
  /* TG68KdotC_Kernel.vhd:671:46  */
  assign n452_o = {1'b0, n450_o};
  /* TG68KdotC_Kernel.vhd:673:53  */
  assign n453_o = sndopc[14:12];
  /* TG68KdotC_Kernel.vhd:673:46  */
  assign n455_o = {1'b0, n453_o};
  /* TG68KdotC_Kernel.vhd:675:53  */
  assign n456_o = sndopc[8:6];
  /* TG68KdotC_Kernel.vhd:675:46  */
  assign n458_o = {1'b0, n456_o};
  /* TG68KdotC_Kernel.vhd:677:61  */
  assign n459_o = last_data_read[2:0];
  /* TG68KdotC_Kernel.vhd:677:46  */
  assign n461_o = {1'b0, n459_o};
  /* TG68KdotC_Kernel.vhd:679:61  */
  assign n462_o = last_data_read[8:6];
  /* TG68KdotC_Kernel.vhd:679:46  */
  assign n464_o = {1'b0, n462_o};
  /* TG68KdotC_Kernel.vhd:681:61  */
  assign n465_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:681:54  */
  assign n466_o = {source_areg, n465_o};
  /* TG68KdotC_Kernel.vhd:682:27  */
  assign n467_o = exec[36];
  /* TG68KdotC_Kernel.vhd:685:61  */
  assign n468_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:685:54  */
  assign n469_o = {source_areg, n468_o};
  /* TG68KdotC_Kernel.vhd:682:17  */
  assign n471_o = n467_o ? 4'b1111 : n469_o;
  /* TG68KdotC_Kernel.vhd:680:17  */
  assign n472_o = source_lowbits ? n466_o : n471_o;
  /* TG68KdotC_Kernel.vhd:678:17  */
  assign n473_o = source_ldrmbits ? n464_o : n472_o;
  /* TG68KdotC_Kernel.vhd:676:17  */
  assign n474_o = source_ldrlbits ? n461_o : n473_o;
  /* TG68KdotC_Kernel.vhd:674:17  */
  assign n475_o = source_2ndmbits ? n458_o : n474_o;
  /* TG68KdotC_Kernel.vhd:672:17  */
  assign n476_o = source_2ndhbits ? n455_o : n475_o;
  /* TG68KdotC_Kernel.vhd:670:17  */
  assign n477_o = source_2ndlbits ? n452_o : n476_o;
  /* TG68KdotC_Kernel.vhd:664:17  */
  assign n478_o = n446_o ? n449_o : n477_o;
  /* TG68KdotC_Kernel.vhd:695:24  */
  assign n482_o = exec[54];
  /* TG68KdotC_Kernel.vhd:697:27  */
  assign n483_o = exec[26];
  /* TG68KdotC_Kernel.vhd:697:45  */
  assign n484_o = store_in_tmp & n483_o;
  /* TG68KdotC_Kernel.vhd:699:27  */
  assign n485_o = exec[69];
  /* TG68KdotC_Kernel.vhd:699:59  */
  assign n486_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:699:62  */
  assign n487_o = ~n486_o;
  /* TG68KdotC_Kernel.vhd:699:46  */
  assign n488_o = n485_o | n487_o;
  /* TG68KdotC_Kernel.vhd:699:74  */
  assign n489_o = exec[39];
  /* TG68KdotC_Kernel.vhd:699:67  */
  assign n490_o = n488_o | n489_o;
  /* TG68KdotC_Kernel.vhd:699:17  */
  assign n491_o = n490_o ? addr : reg_qa;
  /* TG68KdotC_Kernel.vhd:697:17  */
  assign n492_o = n484_o ? ea_data : n491_o;
  /* TG68KdotC_Kernel.vhd:695:17  */
  assign n494_o = n482_o ? 32'b00000000000000000000000000000000 : n492_o;
  /* TG68KdotC_Kernel.vhd:710:46  */
  assign n498_o = reg_qb[15:0];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n499_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n500_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n501_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n502_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n503_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n504_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n505_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n506_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n507_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n508_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n509_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n510_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n511_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n512_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n513_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n514_o = op2out[15];
  assign n515_o = {n499_o, n500_o, n501_o, n502_o};
  assign n516_o = {n503_o, n504_o, n505_o, n506_o};
  assign n517_o = {n507_o, n508_o, n509_o, n510_o};
  assign n518_o = {n511_o, n512_o, n513_o, n514_o};
  assign n519_o = {n515_o, n516_o, n517_o, n518_o};
  /* TG68KdotC_Kernel.vhd:712:24  */
  assign n520_o = exec[53];
  /* TG68KdotC_Kernel.vhd:714:51  */
  assign n522_o = exec[61];
  /* TG68KdotC_Kernel.vhd:714:61  */
  assign n523_o = execopc & n522_o;
  /* TG68KdotC_Kernel.vhd:714:43  */
  assign n524_o = use_direct_data | n523_o;
  /* TG68KdotC_Kernel.vhd:714:85  */
  assign n525_o = exec[29];
  /* TG68KdotC_Kernel.vhd:714:78  */
  assign n526_o = n524_o | n525_o;
  /* TG68KdotC_Kernel.vhd:716:28  */
  assign n527_o = exec[26];
  /* TG68KdotC_Kernel.vhd:716:41  */
  assign n528_o = ~n527_o;
  /* TG68KdotC_Kernel.vhd:716:46  */
  assign n529_o = store_in_tmp & n528_o;
  /* TG68KdotC_Kernel.vhd:716:75  */
  assign n530_o = exec[27];
  /* TG68KdotC_Kernel.vhd:716:68  */
  assign n531_o = n529_o | n530_o;
  /* TG68KdotC_Kernel.vhd:718:27  */
  assign n532_o = exec[1];
  /* TG68KdotC_Kernel.vhd:719:57  */
  assign n533_o = exe_opcode[7:0];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n534_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n535_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n536_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n537_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n538_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n539_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n540_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n541_o = exe_opcode[7];
  assign n542_o = {n534_o, n535_o, n536_o, n537_o};
  assign n543_o = {n538_o, n539_o, n540_o, n541_o};
  assign n544_o = {n542_o, n543_o};
  /* TG68KdotC_Kernel.vhd:721:27  */
  assign n545_o = exec[4];
  /* TG68KdotC_Kernel.vhd:722:57  */
  assign n546_o = exe_opcode[11:9];
  /* TG68KdotC_Kernel.vhd:723:38  */
  assign n547_o = exe_opcode[11:9];
  /* TG68KdotC_Kernel.vhd:723:51  */
  assign n549_o = n547_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:723:25  */
  assign n552_o = n549_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:729:35  */
  assign n555_o = exe_datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:729:49  */
  assign n556_o = exec[11];
  /* TG68KdotC_Kernel.vhd:729:57  */
  assign n557_o = ~n556_o;
  /* TG68KdotC_Kernel.vhd:729:41  */
  assign n558_o = n557_o & n555_o;
  /* TG68KdotC_Kernel.vhd:730:55  */
  assign n559_o = reg_qb[31:16];
  /* TG68KdotC_Kernel.vhd:729:17  */
  assign n560_o = n558_o ? n559_o : n519_o;
  assign n561_o = {12'b000000000000, n552_o, n546_o};
  /* TG68KdotC_Kernel.vhd:721:17  */
  assign n562_o = n545_o ? n561_o : n498_o;
  /* TG68KdotC_Kernel.vhd:721:17  */
  assign n563_o = n545_o ? n519_o : n560_o;
  assign n564_o = {n563_o, n562_o};
  assign n565_o = {n544_o, n533_o};
  assign n566_o = n564_o[15:0];
  /* TG68KdotC_Kernel.vhd:718:17  */
  assign n567_o = n532_o ? n565_o : n566_o;
  assign n568_o = n564_o[31:16];
  /* TG68KdotC_Kernel.vhd:718:17  */
  assign n569_o = n532_o ? n519_o : n568_o;
  assign n570_o = {n569_o, n567_o};
  /* TG68KdotC_Kernel.vhd:716:17  */
  assign n571_o = n531_o ? ea_data : n570_o;
  /* TG68KdotC_Kernel.vhd:714:17  */
  assign n572_o = n526_o ? data_write_tmp : n571_o;
  assign n575_o = n572_o[31:16];
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n576_o = n520_o ? n519_o : n575_o;
  /* TG68KdotC_Kernel.vhd:732:24  */
  assign n577_o = exec[88];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n578_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n579_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n580_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n581_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n582_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n583_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n584_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n585_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n586_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n587_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n588_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n589_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n590_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n591_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n592_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n593_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n594_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n595_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n596_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n597_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n598_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n599_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n600_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n601_o = op2out[7];
  assign n602_o = {n578_o, n579_o, n580_o, n581_o};
  assign n603_o = {n582_o, n583_o, n584_o, n585_o};
  assign n604_o = {n586_o, n587_o, n588_o, n589_o};
  assign n605_o = {n590_o, n591_o, n592_o, n593_o};
  assign n606_o = {n594_o, n595_o, n596_o, n597_o};
  assign n607_o = {n598_o, n599_o, n600_o, n601_o};
  assign n608_o = {n602_o, n603_o, n604_o, n605_o};
  assign n609_o = {n606_o, n607_o};
  assign n610_o = {n608_o, n609_o};
  assign n611_o = n521_o[15:8];
  assign n612_o = data_write_tmp[15:8];
  assign n613_o = ea_data[15:8];
  assign n614_o = n570_o[15:8];
  /* TG68KdotC_Kernel.vhd:716:17  */
  assign n615_o = n531_o ? n613_o : n614_o;
  /* TG68KdotC_Kernel.vhd:714:17  */
  assign n616_o = n526_o ? n612_o : n615_o;
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n617_o = n520_o ? n611_o : n616_o;
  assign n618_o = {n576_o, n617_o};
  /* TG68KdotC_Kernel.vhd:732:17  */
  assign n619_o = n577_o ? n610_o : n618_o;
  assign n620_o = n521_o[7:0];
  assign n621_o = data_write_tmp[7:0];
  assign n622_o = ea_data[7:0];
  assign n623_o = n570_o[7:0];
  /* TG68KdotC_Kernel.vhd:716:17  */
  assign n624_o = n531_o ? n622_o : n623_o;
  /* TG68KdotC_Kernel.vhd:714:17  */
  assign n625_o = n526_o ? n621_o : n624_o;
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n626_o = n520_o ? n620_o : n625_o;
  /* TG68KdotC_Kernel.vhd:753:40  */
  assign n631_o = exec[82];
  /* TG68KdotC_Kernel.vhd:753:33  */
  assign n633_o = n631_o ? 1'b1 : use_direct_data;
  /* TG68KdotC_Kernel.vhd:759:56  */
  assign n634_o = set[27];
  /* TG68KdotC_Kernel.vhd:759:50  */
  assign n635_o = endopc | n634_o;
  /* TG68KdotC_Kernel.vhd:759:33  */
  assign n637_o = n635_o ? 1'b0 : n633_o;
  /* TG68KdotC_Kernel.vhd:756:33  */
  assign n639_o = set_direct_data ? 1'b1 : n637_o;
  /* TG68KdotC_Kernel.vhd:756:33  */
  assign n642_o = set_direct_data ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:762:56  */
  assign n644_o = set_exec[0];
  /* TG68KdotC_Kernel.vhd:769:41  */
  assign n646_o = set_z_error ? 1'b1 : z_error;
  /* TG68KdotC_Kernel.vhd:772:52  */
  assign n647_o = set_exec[0];
  /* TG68KdotC_Kernel.vhd:772:75  */
  assign n649_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:772:66  */
  assign n650_o = n649_o & n647_o;
  /* TG68KdotC_Kernel.vhd:772:41  */
  assign n652_o = n650_o ? 1'b1 : n639_o;
  /* TG68KdotC_Kernel.vhd:776:49  */
  assign n654_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:776:62  */
  assign n655_o = exec[80];
  /* TG68KdotC_Kernel.vhd:776:55  */
  assign n656_o = n654_o | n655_o;
  /* TG68KdotC_Kernel.vhd:776:41  */
  assign n658_o = n656_o ? 1'b1 : store_in_tmp;
  /* TG68KdotC_Kernel.vhd:779:69  */
  assign n660_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:779:60  */
  assign n661_o = n660_o & direct_data;
  /* TG68KdotC_Kernel.vhd:779:41  */
  assign n663_o = n661_o ? 1'b1 : n658_o;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n665_o = endopc ? 1'b0 : n663_o;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n667_o = endopc ? 1'b0 : writepcnext;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n668_o = endopc ? n639_o : n652_o;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n670_o = endopc ? 1'b0 : n646_o;
  /* TG68KdotC_Kernel.vhd:784:41  */
  assign n672_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:784:55  */
  assign n673_o = exec[79];
  /* TG68KdotC_Kernel.vhd:784:69  */
  assign n674_o = ~n673_o;
  /* TG68KdotC_Kernel.vhd:784:47  */
  assign n675_o = n674_o & n672_o;
  /* TG68KdotC_Kernel.vhd:786:43  */
  assign n676_o = exec[71];
  /* TG68KdotC_Kernel.vhd:788:43  */
  assign n677_o = exec[44];
  /* TG68KdotC_Kernel.vhd:788:92  */
  assign n679_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:788:83  */
  assign n680_o = n679_o & direct_data;
  /* TG68KdotC_Kernel.vhd:788:63  */
  assign n681_o = n677_o | n680_o;
  /* TG68KdotC_Kernel.vhd:788:33  */
  assign n682_o = n681_o ? last_data_read : ea_data;
  /* TG68KdotC_Kernel.vhd:786:33  */
  assign n683_o = n676_o ? addr : n682_o;
  /* TG68KdotC_Kernel.vhd:784:33  */
  assign n684_o = n675_o ? data_read : n683_o;
  /* TG68KdotC_Kernel.vhd:794:43  */
  assign n685_o = exec[25];
  /* TG68KdotC_Kernel.vhd:797:50  */
  assign n687_o = $unsigned(micro_state) >= $unsigned(7'b1000110);
  /* TG68KdotC_Kernel.vhd:797:74  */
  assign n689_o = $unsigned(micro_state) <= $unsigned(7'b1011110);
  /* TG68KdotC_Kernel.vhd:797:58  */
  assign n690_o = n689_o & n687_o;
  /* TG68KdotC_Kernel.vhd:799:50  */
  assign n692_o = micro_state == 7'b0110010;
  /* TG68KdotC_Kernel.vhd:802:66  */
  assign n693_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:802:87  */
  assign n694_o = exec[43];
  /* TG68KdotC_Kernel.vhd:802:80  */
  assign n695_o = n693_o | n694_o;
  /* TG68KdotC_Kernel.vhd:802:98  */
  assign n696_o = n695_o | z_error;
  /* TG68KdotC_Kernel.vhd:803:51  */
  assign n698_o = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:809:100  */
  assign n699_o = trap_vector[11:0];
  /* TG68KdotC_Kernel.vhd:809:87  */
  assign n701_o = {4'b0010, n699_o};
  /* TG68KdotC_Kernel.vhd:811:61  */
  assign n702_o = trap_berr | trap_addr_error;
  /* TG68KdotC_Kernel.vhd:812:100  */
  assign n703_o = trap_vector[11:0];
  /* TG68KdotC_Kernel.vhd:812:87  */
  assign n705_o = {4'b1111, n703_o};
  /* TG68KdotC_Kernel.vhd:813:74  */
  assign n706_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:813:95  */
  assign n707_o = exec[43];
  /* TG68KdotC_Kernel.vhd:813:88  */
  assign n708_o = n706_o | n707_o;
  /* TG68KdotC_Kernel.vhd:813:106  */
  assign n709_o = n708_o | z_error;
  /* TG68KdotC_Kernel.vhd:815:100  */
  assign n710_o = trap_vector[11:0];
  /* TG68KdotC_Kernel.vhd:815:87  */
  assign n712_o = {4'b0000, n710_o};
  /* TG68KdotC_Kernel.vhd:816:74  */
  assign n713_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:816:95  */
  assign n714_o = exec[43];
  /* TG68KdotC_Kernel.vhd:816:88  */
  assign n715_o = n713_o | n714_o;
  /* TG68KdotC_Kernel.vhd:816:106  */
  assign n716_o = n715_o | z_error;
  /* TG68KdotC_Kernel.vhd:811:41  */
  assign n717_o = n702_o ? n705_o : n712_o;
  /* TG68KdotC_Kernel.vhd:811:41  */
  assign n718_o = n702_o ? n709_o : n716_o;
  /* TG68KdotC_Kernel.vhd:807:41  */
  assign n719_o = usestackframe2 ? n701_o : n717_o;
  /* TG68KdotC_Kernel.vhd:807:41  */
  assign n720_o = usestackframe2 ? n667_o : n718_o;
  /* TG68KdotC_Kernel.vhd:821:43  */
  assign n721_o = exec[64];
  /* TG68KdotC_Kernel.vhd:823:43  */
  assign n722_o = exec[61];
  /* TG68KdotC_Kernel.vhd:825:43  */
  assign n723_o = exec[62];
  /* TG68KdotC_Kernel.vhd:825:60  */
  assign n724_o = ea_only & n723_o;
  /* TG68KdotC_Kernel.vhd:829:65  */
  assign n726_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:829:56  */
  assign n727_o = n726_o & exec_direct;
  /* TG68KdotC_Kernel.vhd:831:49  */
  assign n728_o = exec[37];
  /* TG68KdotC_Kernel.vhd:832:94  */
  assign n729_o = data_write_tmp[23:0];
  assign n730_o = data_read[31:8];
  /* TG68KdotC_Kernel.vhd:831:41  */
  assign n731_o = n728_o ? n729_o : n730_o;
  assign n732_o = data_read[7:0];
  /* TG68KdotC_Kernel.vhd:834:43  */
  assign n733_o = exec[37];
  /* TG68KdotC_Kernel.vhd:835:78  */
  assign n734_o = reg_qb[31:16];
  /* TG68KdotC_Kernel.vhd:839:91  */
  assign n735_o = {trap_sr, flags};
  assign n736_o = op2out[15:0];
  /* TG68KdotC_Kernel.vhd:838:33  */
  assign n737_o = writesr ? n735_o : n736_o;
  assign n738_o = op2out[31:16];
  assign n739_o = data_write_tmp[31:16];
  /* TG68KdotC_Kernel.vhd:838:33  */
  assign n740_o = writesr ? n739_o : n738_o;
  assign n741_o = {n740_o, n737_o};
  /* TG68KdotC_Kernel.vhd:836:33  */
  assign n742_o = direct_data ? last_data_read : n741_o;
  assign n743_o = n742_o[15:0];
  /* TG68KdotC_Kernel.vhd:834:33  */
  assign n744_o = n733_o ? n734_o : n743_o;
  assign n745_o = n742_o[31:16];
  assign n746_o = data_write_tmp[31:16];
  /* TG68KdotC_Kernel.vhd:834:33  */
  assign n747_o = n733_o ? n746_o : n745_o;
  assign n748_o = {n747_o, n744_o};
  assign n749_o = {n731_o, n732_o};
  /* TG68KdotC_Kernel.vhd:829:33  */
  assign n750_o = n727_o ? n749_o : n748_o;
  /* TG68KdotC_Kernel.vhd:827:33  */
  assign n751_o = execopc ? aluout : n750_o;
  /* TG68KdotC_Kernel.vhd:825:33  */
  assign n752_o = n724_o ? addr : n751_o;
  /* TG68KdotC_Kernel.vhd:823:33  */
  assign n753_o = n722_o ? op1out : n752_o;
  /* TG68KdotC_Kernel.vhd:821:33  */
  assign n754_o = n721_o ? data_write_tmp : n753_o;
  assign n755_o = n754_o[15:0];
  /* TG68KdotC_Kernel.vhd:803:33  */
  assign n756_o = n698_o ? n719_o : n755_o;
  assign n757_o = n754_o[31:16];
  assign n758_o = data_write_tmp[31:16];
  /* TG68KdotC_Kernel.vhd:803:33  */
  assign n759_o = n698_o ? n758_o : n757_o;
  /* TG68KdotC_Kernel.vhd:803:33  */
  assign n760_o = n698_o ? n720_o : n667_o;
  assign n761_o = {n759_o, n756_o};
  /* TG68KdotC_Kernel.vhd:799:33  */
  assign n762_o = n692_o ? exe_pc : n761_o;
  /* TG68KdotC_Kernel.vhd:799:33  */
  assign n763_o = n692_o ? n696_o : n760_o;
  /* TG68KdotC_Kernel.vhd:799:33  */
  assign n766_o = n692_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n768_o = n690_o ? 32'b00000000000000000000000000000000 : n762_o;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n769_o = n690_o ? n667_o : n763_o;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n771_o = n690_o ? 1'b0 : n766_o;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n772_o = n685_o ? tg68_pc_add : n768_o;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n773_o = n685_o ? n667_o : n769_o;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n775_o = n685_o ? 1'b0 : n771_o;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n776_o = writepc ? tg68_pc : n772_o;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n777_o = writepc ? n667_o : n773_o;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n779_o = writepc ? 1'b0 : n775_o;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n781_o = clkena_lw ? n684_o : ea_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n782_o = clkena_lw ? n776_o : data_write_tmp;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n783_o = clkena_lw ? n665_o : store_in_tmp;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n784_o = clkena_lw ? n777_o : writepcnext;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n785_o = clkena_lw ? n644_o : exec_direct;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n786_o = clkena_lw ? n668_o : use_direct_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n787_o = clkena_lw ? n642_o : direct_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n788_o = clkena_lw ? n779_o : usestackframe2;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n789_o = clkena_lw ? n670_o : z_error;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n790_o = reset ? ea_data : n781_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n791_o = reset ? data_write_tmp : n782_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n793_o = reset ? 1'b0 : n783_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n795_o = reset ? 1'b0 : n784_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n796_o = reset ? exec_direct : n785_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n798_o = reset ? 1'b0 : n786_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n800_o = reset ? 1'b0 : n787_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n801_o = reset ? usestackframe2 : n788_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n803_o = reset ? 1'b0 : n789_o;
  /* TG68KdotC_Kernel.vhd:852:25  */
  assign n816_o = brief[11];
  /* TG68KdotC_Kernel.vhd:853:46  */
  assign n817_o = op1out[31:16];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n818_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n819_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n820_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n821_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n822_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n823_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n824_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n825_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n826_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n827_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n828_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n829_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n830_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n831_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n832_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n833_o = op1out[15];
  assign n834_o = {n818_o, n819_o, n820_o, n821_o};
  assign n835_o = {n822_o, n823_o, n824_o, n825_o};
  assign n836_o = {n826_o, n827_o, n828_o, n829_o};
  assign n837_o = {n830_o, n831_o, n832_o, n833_o};
  assign n838_o = {n834_o, n835_o, n836_o, n837_o};
  /* TG68KdotC_Kernel.vhd:852:17  */
  assign n839_o = n816_o ? n817_o : n838_o;
  /* TG68KdotC_Kernel.vhd:857:48  */
  assign n840_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:857:41  */
  assign n841_o = {op1outbrief, n840_o};
  /* TG68KdotC_Kernel.vhd:858:42  */
  assign n842_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:858:50  */
  assign n844_o = 1'b1 & n842_o;
  /* TG68KdotC_Kernel.vhd:858:35  */
  assign n846_o = 1'b0 | n844_o;
  /* TG68KdotC_Kernel.vhd:859:35  */
  assign n847_o = brief[10:9];
  /* TG68KdotC_Kernel.vhd:860:77  */
  assign n848_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:860:70  */
  assign n849_o = {op1outbrief, n848_o};
  /* TG68KdotC_Kernel.vhd:860:33  */
  assign n851_o = n847_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:861:70  */
  assign n852_o = op1outbrief[14:0];
  /* TG68KdotC_Kernel.vhd:861:90  */
  assign n853_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:861:83  */
  assign n854_o = {n852_o, n853_o};
  /* TG68KdotC_Kernel.vhd:861:103  */
  assign n856_o = {n854_o, 1'b0};
  /* TG68KdotC_Kernel.vhd:861:33  */
  assign n858_o = n847_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:862:70  */
  assign n859_o = op1outbrief[13:0];
  /* TG68KdotC_Kernel.vhd:862:90  */
  assign n860_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:862:83  */
  assign n861_o = {n859_o, n860_o};
  /* TG68KdotC_Kernel.vhd:862:103  */
  assign n863_o = {n861_o, 2'b00};
  /* TG68KdotC_Kernel.vhd:862:33  */
  assign n865_o = n847_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:863:70  */
  assign n866_o = op1outbrief[12:0];
  /* TG68KdotC_Kernel.vhd:863:90  */
  assign n867_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:863:83  */
  assign n868_o = {n866_o, n867_o};
  /* TG68KdotC_Kernel.vhd:863:103  */
  assign n870_o = {n868_o, 3'b000};
  /* TG68KdotC_Kernel.vhd:863:33  */
  assign n872_o = n847_o == 2'b11;
  assign n873_o = {n872_o, n865_o, n858_o, n851_o};
  /* TG68KdotC_Kernel.vhd:859:25  */
  always @*
    case (n873_o)
      4'b1000: n874_o = n870_o;
      4'b0100: n874_o = n863_o;
      4'b0010: n874_o = n856_o;
      4'b0001: n874_o = n849_o;
      default: n874_o = n841_o;
    endcase
  /* TG68KdotC_Kernel.vhd:858:17  */
  assign n875_o = n846_o ? n874_o : n841_o;
  assign n882_o = trap_vector[9:0];
  /* TG68KdotC_Kernel.vhd:879:33  */
  assign n883_o = trap_berr ? 10'b0000001000 : n882_o;
  /* TG68KdotC_Kernel.vhd:882:33  */
  assign n885_o = trap_addr_error ? 10'b0000001100 : n883_o;
  /* TG68KdotC_Kernel.vhd:885:33  */
  assign n887_o = trap_illegal ? 10'b0000010000 : n885_o;
  /* TG68KdotC_Kernel.vhd:888:33  */
  assign n889_o = set_z_error ? 10'b0000010100 : n887_o;
  /* TG68KdotC_Kernel.vhd:891:40  */
  assign n890_o = exec[43];
  /* TG68KdotC_Kernel.vhd:891:33  */
  assign n892_o = n890_o ? 10'b0000011000 : n889_o;
  /* TG68KdotC_Kernel.vhd:894:33  */
  assign n894_o = trap_trapv ? 10'b0000011100 : n892_o;
  /* TG68KdotC_Kernel.vhd:897:33  */
  assign n896_o = trap_priv ? 10'b0000100000 : n894_o;
  /* TG68KdotC_Kernel.vhd:900:33  */
  assign n898_o = trap_trace ? 10'b0000100100 : n896_o;
  /* TG68KdotC_Kernel.vhd:903:33  */
  assign n900_o = trap_1010 ? 10'b0000101000 : n898_o;
  /* TG68KdotC_Kernel.vhd:906:33  */
  assign n902_o = trap_1111 ? 10'b0000101100 : n900_o;
  /* TG68KdotC_Kernel.vhd:910:83  */
  assign n903_o = opcode[3:0];
  /* TG68KdotC_Kernel.vhd:910:75  */
  assign n905_o = {4'b0010, n903_o};
  /* TG68KdotC_Kernel.vhd:910:96  */
  assign n907_o = {n905_o, 2'b00};
  /* TG68KdotC_Kernel.vhd:909:33  */
  assign n908_o = trap_trap ? n907_o : n902_o;
  /* TG68KdotC_Kernel.vhd:912:55  */
  assign n909_o = trap_interrupt | set_vectoraddr;
  /* TG68KdotC_Kernel.vhd:913:76  */
  assign n911_o = {ipl_vec, 2'b00};
  /* TG68KdotC_Kernel.vhd:912:33  */
  assign n912_o = n909_o ? n911_o : n908_o;
  assign n913_o = {22'b0000000000000000000000, n912_o};
  /* TG68KdotC_Kernel.vhd:918:55  */
  assign n916_o = trap_vector + vbr;
  /* TG68KdotC_Kernel.vhd:917:17  */
  assign n917_o = use_vbr_stackframe ? n916_o : trap_vector;
  /* TG68KdotC_Kernel.vhd:924:60  */
  assign n919_o = memaddr_a[4];
  /* TG68KdotC_Kernel.vhd:924:60  */
  assign n920_o = memaddr_a[4];
  /* TG68KdotC_Kernel.vhd:924:60  */
  assign n921_o = memaddr_a[4];
  assign n922_o = {n919_o, n920_o, n921_o};
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n923_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n924_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n925_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n926_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n927_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n928_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n929_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n930_o = memaddr_a[7];
  assign n931_o = {n923_o, n924_o, n925_o, n926_o};
  assign n932_o = {n927_o, n928_o, n929_o, n930_o};
  assign n933_o = {n931_o, n932_o};
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n934_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n935_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n936_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n937_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n938_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n939_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n940_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n941_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n942_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n943_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n944_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n945_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n946_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n947_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n948_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n949_o = memaddr_a[15];
  assign n950_o = {n934_o, n935_o, n936_o, n937_o};
  assign n951_o = {n938_o, n939_o, n940_o, n941_o};
  assign n952_o = {n942_o, n943_o, n944_o, n945_o};
  assign n953_o = {n946_o, n947_o, n948_o, n949_o};
  assign n954_o = {n950_o, n951_o, n952_o, n953_o};
  /* TG68KdotC_Kernel.vhd:928:32  */
  assign n955_o = exec[70];
  /* TG68KdotC_Kernel.vhd:929:55  */
  assign n956_o = briefdata + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:931:72  */
  assign n957_o = last_data_read[7:0];
  assign n958_o = last_data_read[7:0];
  /* TG68KdotC_Kernel.vhd:930:25  */
  assign n959_o = setdispbyte ? n957_o : n958_o;
  assign n960_o = last_data_read[31:8];
  assign n961_o = {n954_o, n933_o};
  /* TG68KdotC_Kernel.vhd:930:25  */
  assign n962_o = setdispbyte ? n961_o : n960_o;
  assign n963_o = {n962_o, n959_o};
  /* TG68KdotC_Kernel.vhd:928:25  */
  assign n964_o = n955_o ? n956_o : n963_o;
  /* TG68KdotC_Kernel.vhd:935:26  */
  assign n965_o = set[47];
  /* TG68KdotC_Kernel.vhd:936:31  */
  assign n966_o = set[73];
  /* TG68KdotC_Kernel.vhd:938:39  */
  assign n969_o = datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:938:52  */
  assign n970_o = set[50];
  /* TG68KdotC_Kernel.vhd:938:60  */
  assign n971_o = ~n970_o;
  /* TG68KdotC_Kernel.vhd:938:45  */
  assign n972_o = n971_o & n969_o;
  /* TG68KdotC_Kernel.vhd:938:25  */
  assign n975_o = n972_o ? 5'b11111 : 5'b11110;
  /* TG68KdotC_Kernel.vhd:936:25  */
  assign n976_o = n966_o ? 5'b11100 : n975_o;
  /* TG68KdotC_Kernel.vhd:944:53  */
  assign n978_o = {1'b1, ripl_nr};
  /* TG68KdotC_Kernel.vhd:944:61  */
  assign n980_o = {n978_o, 1'b0};
  /* TG68KdotC_Kernel.vhd:943:17  */
  assign n981_o = interrupt ? n980_o : 5'b00000;
  /* TG68KdotC_Kernel.vhd:935:17  */
  assign n982_o = n965_o ? n976_o : n981_o;
  assign n983_o = n964_o[4:0];
  /* TG68KdotC_Kernel.vhd:927:17  */
  assign n984_o = setdisp ? n983_o : n982_o;
  assign n985_o = n964_o[31:5];
  assign n986_o = {n954_o, n933_o, n922_o};
  /* TG68KdotC_Kernel.vhd:927:17  */
  assign n987_o = setdisp ? n985_o : n986_o;
  /* TG68KdotC_Kernel.vhd:949:40  */
  assign n989_o = exec[71];
  /* TG68KdotC_Kernel.vhd:949:66  */
  assign n991_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:949:83  */
  assign n992_o = memread[0];
  /* TG68KdotC_Kernel.vhd:949:72  */
  assign n993_o = n992_o & n991_o;
  /* TG68KdotC_Kernel.vhd:949:57  */
  assign n994_o = n989_o | n993_o;
  /* TG68KdotC_Kernel.vhd:954:46  */
  assign n996_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:954:49  */
  assign n997_o = ~n996_o;
  /* TG68KdotC_Kernel.vhd:954:61  */
  assign n998_o = exec[55];
  /* TG68KdotC_Kernel.vhd:954:54  */
  assign n999_o = n997_o | n998_o;
  /* TG68KdotC_Kernel.vhd:956:42  */
  assign n1000_o = set[83];
  /* TG68KdotC_Kernel.vhd:958:43  */
  assign n1001_o = exec[58];
  /* TG68KdotC_Kernel.vhd:960:43  */
  assign n1002_o = exec[63];
  /* TG68KdotC_Kernel.vhd:960:70  */
  assign n1004_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:960:58  */
  assign n1005_o = n1004_o & n1002_o;
  /* TG68KdotC_Kernel.vhd:962:42  */
  assign n1006_o = set[45];
  /* TG68KdotC_Kernel.vhd:964:47  */
  assign n1008_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:966:43  */
  assign n1009_o = exec[22];
  /* TG68KdotC_Kernel.vhd:973:53  */
  assign n1010_o = ~interrupt;
  /* TG68KdotC_Kernel.vhd:973:75  */
  assign n1011_o = ~suppress_base;
  /* TG68KdotC_Kernel.vhd:973:58  */
  assign n1012_o = n1011_o & n1010_o;
  /* TG68KdotC_Kernel.vhd:973:41  */
  assign n1015_o = n1012_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:969:33  */
  assign n1016_o = set_vectoraddr ? trap_vector_vbr : memaddr_a;
  /* TG68KdotC_Kernel.vhd:969:33  */
  assign n1018_o = set_vectoraddr ? 1'b0 : n1015_o;
  /* TG68KdotC_Kernel.vhd:966:33  */
  assign n1019_o = n1009_o ? ea_data : n1016_o;
  /* TG68KdotC_Kernel.vhd:966:33  */
  assign n1021_o = n1009_o ? memaddr_a : 32'b00000000000000000000000000000000;
  /* TG68KdotC_Kernel.vhd:966:33  */
  assign n1023_o = n1009_o ? 1'b0 : n1018_o;
  /* TG68KdotC_Kernel.vhd:964:33  */
  assign n1024_o = n1008_o ? tg68_pc_add : n1019_o;
  /* TG68KdotC_Kernel.vhd:964:33  */
  assign n1026_o = n1008_o ? 32'b00000000000000000000000000000000 : n1021_o;
  /* TG68KdotC_Kernel.vhd:964:33  */
  assign n1028_o = n1008_o ? 1'b0 : n1023_o;
  /* TG68KdotC_Kernel.vhd:962:33  */
  assign n1029_o = n1006_o ? last_data_read : n1024_o;
  /* TG68KdotC_Kernel.vhd:962:33  */
  assign n1031_o = n1006_o ? 32'b00000000000000000000000000000000 : n1026_o;
  /* TG68KdotC_Kernel.vhd:962:33  */
  assign n1033_o = n1006_o ? 1'b0 : n1028_o;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n1034_o = n1005_o ? addr : n1029_o;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n1036_o = n1005_o ? 32'b00000000000000000000000000000000 : n1031_o;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n1038_o = n1005_o ? 1'b0 : n1033_o;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n1039_o = n1001_o ? data_read : n1034_o;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n1041_o = n1001_o ? 32'b00000000000000000000000000000000 : n1036_o;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n1043_o = n1001_o ? 1'b0 : n1038_o;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n1044_o = n1000_o ? tmp_tg68_pc : n1039_o;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n1046_o = n1000_o ? 32'b00000000000000000000000000000000 : n1041_o;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n1048_o = n1000_o ? 1'b0 : n1043_o;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n1049_o = n999_o ? addsub_q : n1044_o;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n1051_o = n999_o ? 32'b00000000000000000000000000000000 : n1046_o;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n1054_o = n999_o ? 1'b0 : n1048_o;
  /* TG68KdotC_Kernel.vhd:981:53  */
  assign n1056_o = memread[0];
  /* TG68KdotC_Kernel.vhd:981:73  */
  assign n1057_o = state[1];
  /* TG68KdotC_Kernel.vhd:981:64  */
  assign n1058_o = n1057_o & n1056_o;
  /* TG68KdotC_Kernel.vhd:981:100  */
  assign n1059_o = ~movem_presub;
  /* TG68KdotC_Kernel.vhd:981:84  */
  assign n1060_o = n1058_o | n1059_o;
  /* TG68KdotC_Kernel.vhd:948:25  */
  assign n1062_o = n994_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:948:25  */
  assign n1063_o = n1060_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:987:53  */
  assign n1072_o = memaddr_delta_rega + memaddr_delta_regb;
  /* TG68KdotC_Kernel.vhd:989:36  */
  assign n1073_o = memaddr_reg + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:990:41  */
  assign n1074_o = memaddr_reg + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:992:28  */
  assign n1075_o = ~use_base;
  /* TG68KdotC_Kernel.vhd:992:17  */
  assign n1077_o = n1075_o ? 32'b00000000000000000000000000000000 : reg_qa;
  /* TG68KdotC_Kernel.vhd:1007:17  */
  assign n1081_o = tg68_pc_brw ? tmp_tg68_pc : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1012:40  */
  assign n1083_o = pc_datab[2];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1084_o = pc_datab[3];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1085_o = pc_datab[3];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1086_o = pc_datab[3];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1087_o = pc_datab[3];
  assign n1088_o = {n1084_o, n1085_o, n1086_o, n1087_o};
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1089_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1090_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1091_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1092_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1093_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1094_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1095_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1096_o = pc_datab[7];
  assign n1097_o = {n1089_o, n1090_o, n1091_o, n1092_o};
  assign n1098_o = {n1093_o, n1094_o, n1095_o, n1096_o};
  assign n1099_o = {n1097_o, n1098_o};
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1100_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1101_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1102_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1103_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1104_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1105_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1106_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1107_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1108_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1109_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1110_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1111_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1112_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1113_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1114_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1115_o = pc_datab[15];
  assign n1116_o = {n1100_o, n1101_o, n1102_o, n1103_o};
  assign n1117_o = {n1104_o, n1105_o, n1106_o, n1107_o};
  assign n1118_o = {n1108_o, n1109_o, n1110_o, n1111_o};
  assign n1119_o = {n1112_o, n1113_o, n1114_o, n1115_o};
  assign n1120_o = {n1116_o, n1117_o, n1118_o, n1119_o};
  assign n1124_o = n1082_o[0];
  /* TG68KdotC_Kernel.vhd:1019:24  */
  assign n1125_o = exec[25];
  assign n1129_o = n1121_o[0];
  assign n1130_o = n1082_o[1];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1131_o = interrupt ? n1129_o : n1130_o;
  /* TG68KdotC_Kernel.vhd:1020:25  */
  assign n1132_o = writepcbig ? 1'b1 : n1131_o;
  assign n1133_o = n1121_o[1];
  assign n1134_o = n1082_o[2];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1135_o = interrupt ? n1133_o : n1134_o;
  /* TG68KdotC_Kernel.vhd:1020:25  */
  assign n1136_o = writepcbig ? n1135_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1020:25  */
  assign n1137_o = writepcbig ? 1'b1 : n1083_o;
  /* TG68KdotC_Kernel.vhd:1026:47  */
  assign n1138_o = ~use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:1026:71  */
  assign n1139_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:1026:96  */
  assign n1140_o = exec[43];
  /* TG68KdotC_Kernel.vhd:1026:89  */
  assign n1141_o = n1139_o | n1140_o;
  /* TG68KdotC_Kernel.vhd:1026:111  */
  assign n1142_o = n1141_o | z_error;
  /* TG68KdotC_Kernel.vhd:1026:52  */
  assign n1143_o = n1142_o & n1138_o;
  /* TG68KdotC_Kernel.vhd:1026:128  */
  assign n1144_o = n1143_o | writepcnext;
  /* TG68KdotC_Kernel.vhd:1026:25  */
  assign n1146_o = n1144_o ? 1'b1 : n1132_o;
  /* TG68KdotC_Kernel.vhd:1029:28  */
  assign n1148_o = state == 2'b00;
  assign n1150_o = n1121_o[0];
  assign n1151_o = n1082_o[1];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1152_o = interrupt ? n1150_o : n1151_o;
  /* TG68KdotC_Kernel.vhd:1029:17  */
  assign n1153_o = n1148_o ? 1'b1 : n1152_o;
  assign n1154_o = {n1137_o, n1136_o, n1146_o};
  assign n1155_o = n1154_o[0];
  /* TG68KdotC_Kernel.vhd:1019:17  */
  assign n1156_o = n1125_o ? n1155_o : n1153_o;
  assign n1157_o = n1154_o[2:1];
  assign n1158_o = n1121_o[1];
  assign n1159_o = n1082_o[2];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1160_o = interrupt ? n1158_o : n1159_o;
  assign n1161_o = {n1083_o, n1160_o};
  /* TG68KdotC_Kernel.vhd:1019:17  */
  assign n1162_o = n1125_o ? n1157_o : n1161_o;
  /* TG68KdotC_Kernel.vhd:1036:63  */
  assign n1166_o = opcode[7:0];
  assign n1167_o = last_data_read[7:0];
  /* TG68KdotC_Kernel.vhd:1033:25  */
  assign n1168_o = tg68_pc_word ? n1167_o : n1166_o;
  assign n1169_o = last_data_read[31:8];
  assign n1170_o = {n1120_o, n1099_o};
  /* TG68KdotC_Kernel.vhd:1033:25  */
  assign n1171_o = tg68_pc_word ? n1169_o : n1170_o;
  assign n1172_o = {n1171_o, n1168_o};
  assign n1173_o = {n1120_o, n1099_o, n1088_o, n1162_o, n1156_o, n1124_o};
  /* TG68KdotC_Kernel.vhd:1032:17  */
  assign n1174_o = tg68_pc_brw ? n1172_o : n1173_o;
  /* TG68KdotC_Kernel.vhd:1040:40  */
  assign n1175_o = pc_dataa + pc_datab;
  /* TG68KdotC_Kernel.vhd:1045:28  */
  assign n1177_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1045:54  */
  assign n1179_o = next_micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1045:34  */
  assign n1180_o = n1179_o & n1177_o;
  /* TG68KdotC_Kernel.vhd:1045:75  */
  assign n1181_o = ~setnextpass;
  /* TG68KdotC_Kernel.vhd:1045:60  */
  assign n1182_o = n1181_o & n1180_o;
  /* TG68KdotC_Kernel.vhd:1045:100  */
  assign n1183_o = ~exec_write_back;
  /* TG68KdotC_Kernel.vhd:1045:113  */
  assign n1185_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:1045:105  */
  assign n1186_o = n1183_o | n1185_o;
  /* TG68KdotC_Kernel.vhd:1045:80  */
  assign n1187_o = n1186_o & n1182_o;
  /* TG68KdotC_Kernel.vhd:1045:135  */
  assign n1189_o = set_rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:1045:120  */
  assign n1190_o = n1189_o & n1187_o;
  /* TG68KdotC_Kernel.vhd:1045:157  */
  assign n1191_o = set_exec[31];
  /* TG68KdotC_Kernel.vhd:1045:165  */
  assign n1192_o = ~n1191_o;
  /* TG68KdotC_Kernel.vhd:1045:145  */
  assign n1193_o = n1192_o & n1190_o;
  /* TG68KdotC_Kernel.vhd:1047:35  */
  assign n1194_o = flagssr[2:0];
  /* TG68KdotC_Kernel.vhd:1047:47  */
  assign n1195_o = $unsigned(n1194_o) < $unsigned(ipl_nr);
  /* TG68KdotC_Kernel.vhd:1047:64  */
  assign n1197_o = ipl_nr == 3'b111;
  /* TG68KdotC_Kernel.vhd:1047:55  */
  assign n1198_o = n1195_o | n1197_o;
  /* TG68KdotC_Kernel.vhd:1047:72  */
  assign n1199_o = n1198_o | make_trace;
  /* TG68KdotC_Kernel.vhd:1047:90  */
  assign n1200_o = n1199_o | make_berr;
  /* TG68KdotC_Kernel.vhd:1049:35  */
  assign n1201_o = ~stop;
  /* TG68KdotC_Kernel.vhd:1049:25  */
  assign n1204_o = n1201_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1047:25  */
  assign n1206_o = n1200_o ? 1'b0 : n1204_o;
  /* TG68KdotC_Kernel.vhd:1047:25  */
  assign n1209_o = n1200_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1045:17  */
  assign n1211_o = n1193_o ? n1206_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1045:17  */
  assign n1215_o = n1193_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1045:17  */
  assign n1218_o = n1193_o ? n1209_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1054:28  */
  assign n1221_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1054:54  */
  assign n1223_o = next_micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1054:34  */
  assign n1224_o = n1223_o & n1221_o;
  /* TG68KdotC_Kernel.vhd:1054:79  */
  assign n1225_o = ~set_direct_data;
  /* TG68KdotC_Kernel.vhd:1054:60  */
  assign n1226_o = n1225_o & n1224_o;
  /* TG68KdotC_Kernel.vhd:1054:104  */
  assign n1227_o = ~exec_write_back;
  /* TG68KdotC_Kernel.vhd:1054:118  */
  assign n1229_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1054:137  */
  assign n1230_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:1054:124  */
  assign n1231_o = n1230_o & n1229_o;
  /* TG68KdotC_Kernel.vhd:1054:109  */
  assign n1232_o = n1227_o | n1231_o;
  /* TG68KdotC_Kernel.vhd:1054:84  */
  assign n1233_o = n1232_o & n1226_o;
  /* TG68KdotC_Kernel.vhd:1054:17  */
  assign n1236_o = n1233_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1058:27  */
  assign n1238_o = ~ipl;
  /* TG68KdotC_Kernel.vhd:1088:59  */
  assign n1240_o = memmask[3:0];
  /* TG68KdotC_Kernel.vhd:1088:71  */
  assign n1242_o = {n1240_o, 2'b11};
  /* TG68KdotC_Kernel.vhd:1089:59  */
  assign n1243_o = memread[1:0];
  /* TG68KdotC_Kernel.vhd:1089:82  */
  assign n1244_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:1089:71  */
  assign n1245_o = {n1243_o, n1244_o};
  /* TG68KdotC_Kernel.vhd:1093:48  */
  assign n1246_o = exec[57];
  /* TG68KdotC_Kernel.vhd:1095:51  */
  assign n1247_o = exec[63];
  /* TG68KdotC_Kernel.vhd:1097:54  */
  assign n1249_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1097:60  */
  assign n1250_o = n1249_o | tg68_pc_brw;
  /* TG68KdotC_Kernel.vhd:1097:90  */
  assign n1251_o = ~stop;
  /* TG68KdotC_Kernel.vhd:1097:82  */
  assign n1252_o = n1251_o & n1250_o;
  /* TG68KdotC_Kernel.vhd:1097:41  */
  assign n1253_o = n1252_o ? tg68_pc_add : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1095:41  */
  assign n1254_o = n1247_o ? addr : n1253_o;
  /* TG68KdotC_Kernel.vhd:1093:41  */
  assign n1255_o = n1246_o ? data_read : n1254_o;
  /* TG68KdotC_Kernel.vhd:1087:33  */
  assign n1256_o = clkena_in ? n1255_o : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1087:33  */
  assign n1257_o = clkena_in ? n1242_o : memmask;
  /* TG68KdotC_Kernel.vhd:1087:33  */
  assign n1258_o = clkena_in ? n1245_o : memread;
  /* TG68KdotC_Kernel.vhd:1115:53  */
  assign n1259_o = ~trap_berr;
  /* TG68KdotC_Kernel.vhd:1116:68  */
  assign n1260_o = berr | make_berr;
  /* TG68KdotC_Kernel.vhd:1115:41  */
  assign n1262_o = n1259_o ? n1260_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1121:71  */
  assign n1263_o = ~setinterrupt;
  /* TG68KdotC_Kernel.vhd:1121:67  */
  assign n1264_o = n1263_o & stop;
  /* TG68KdotC_Kernel.vhd:1121:58  */
  assign n1265_o = set_stop | n1264_o;
  /* TG68KdotC_Kernel.vhd:1134:75  */
  assign n1267_o = {5'b00011, ipl_nr};
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1270_o = make_berr ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1273_o = make_berr ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1274_o = make_berr ? ripl_nr : ipl_nr;
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1275_o = make_berr ? ipl_vec : n1267_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1277_o = make_trace ? 1'b0 : n1270_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1281_o = make_trace ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1284_o = make_trace ? 1'b0 : n1273_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1286_o = make_trace ? ripl_nr : n1274_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1287_o = make_trace ? ipl_vec : n1275_o;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1288_o = setinterrupt ? n1277_o : trap_berr;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1289_o = setinterrupt ? n1281_o : trap_trace;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1290_o = setinterrupt ? n1284_o : trap_interrupt;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1292_o = setinterrupt ? 1'b0 : n1262_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1293_o = n1496_o ? n1286_o : ripl_nr;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1294_o = setinterrupt ? n1287_o : ipl_vec;
  /* TG68KdotC_Kernel.vhd:1138:55  */
  assign n1296_o = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1138:80  */
  assign n1297_o = ~ipl_autovector;
  /* TG68KdotC_Kernel.vhd:1138:62  */
  assign n1298_o = n1297_o & n1296_o;
  /* TG68KdotC_Kernel.vhd:1139:74  */
  assign n1299_o = last_data_read[7:0];
  /* TG68KdotC_Kernel.vhd:1138:41  */
  assign n1300_o = n1298_o ? n1299_o : n1294_o;
  /* TG68KdotC_Kernel.vhd:1141:49  */
  assign n1302_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1142:75  */
  assign n1303_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1304_o = n1478_o ? tg68_pc : last_opc_pc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1305_o = n1479_o ? n1303_o : last_opc_read;
  /* TG68KdotC_Kernel.vhd:1150:53  */
  assign n1306_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:1150:65  */
  assign n1308_o = n1306_o == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:1150:86  */
  assign n1309_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:1150:98  */
  assign n1311_o = n1309_o == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:1150:77  */
  assign n1312_o = n1308_o | n1311_o;
  /* TG68KdotC_Kernel.vhd:1150:110  */
  assign n1313_o = n1312_o | data_is_source;
  /* TG68KdotC_Kernel.vhd:1150:41  */
  assign n1315_o = n1313_o ? 1'b1 : tg68_pc_word;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1317_o = setopcode ? 1'b0 : n1315_o;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1319_o = setopcode ? 1'b0 : n1288_o;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1321_o = setopcode ? 1'b0 : n1289_o;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1323_o = setopcode ? 1'b0 : n1290_o;
  /* TG68KdotC_Kernel.vhd:1154:48  */
  assign n1324_o = exec[29];
  /* TG68KdotC_Kernel.vhd:1158:84  */
  assign n1325_o = {26'b0, bf_width};  //  uext
  /* TG68KdotC_Kernel.vhd:1158:84  */
  assign n1326_o = bf_full_offset + n1325_o;
  /* TG68KdotC_Kernel.vhd:1158:93  */
  assign n1328_o = n1326_o + 32'b00000000000000000000000000000001;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1329_o = n1505_o ? bf_width : alu_width;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1330_o = n1506_o ? bf_shift : alu_bf_shift;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1331_o = n1507_o ? n1328_o : alu_bf_ffo_offset;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1332_o = n1508_o ? bf_loffset : alu_bf_loffset;
  /* TG68KdotC_Kernel.vhd:1161:62  */
  assign n1333_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1161:50  */
  assign n1334_o = ~n1333_o;
  /* TG68KdotC_Kernel.vhd:1161:93  */
  assign n1335_o = setstate[0];
  /* TG68KdotC_Kernel.vhd:1161:81  */
  assign n1336_o = ~n1335_o;
  /* TG68KdotC_Kernel.vhd:1161:77  */
  assign n1337_o = pcbase & n1336_o;
  /* TG68KdotC_Kernel.vhd:1161:66  */
  assign n1338_o = n1334_o | n1337_o;
  /* TG68KdotC_Kernel.vhd:1162:58  */
  assign n1339_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1162:67  */
  assign n1340_o = ~pcbase;
  /* TG68KdotC_Kernel.vhd:1162:89  */
  assign n1341_o = setstate[0];
  /* TG68KdotC_Kernel.vhd:1162:78  */
  assign n1342_o = n1340_o | n1341_o;
  /* TG68KdotC_Kernel.vhd:1162:62  */
  assign n1343_o = n1339_o & n1342_o;
  assign n1345_o = {n1338_o, n1343_o};
  /* TG68KdotC_Kernel.vhd:1163:41  */
  assign n1346_o = interrupt ? 2'b11 : n1345_o;
  /* TG68KdotC_Kernel.vhd:1167:49  */
  assign n1348_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:1169:55  */
  assign n1350_o = setstate == 2'b10;
  /* TG68KdotC_Kernel.vhd:1169:77  */
  assign n1351_o = ~setaddrvalue;
  /* TG68KdotC_Kernel.vhd:1169:61  */
  assign n1352_o = n1351_o & n1350_o;
  /* TG68KdotC_Kernel.vhd:1169:82  */
  assign n1353_o = write_back & n1352_o;
  /* TG68KdotC_Kernel.vhd:1169:41  */
  assign n1355_o = n1353_o ? 1'b1 : exec_write_back;
  /* TG68KdotC_Kernel.vhd:1167:41  */
  assign n1357_o = n1348_o ? 1'b0 : n1355_o;
  /* TG68KdotC_Kernel.vhd:1172:50  */
  assign n1359_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1172:69  */
  assign n1360_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:1172:56  */
  assign n1361_o = n1360_o & n1359_o;
  /* TG68KdotC_Kernel.vhd:1172:74  */
  assign n1362_o = write_back & n1361_o;
  /* TG68KdotC_Kernel.vhd:1172:105  */
  assign n1364_o = setstate != 2'b10;
  /* TG68KdotC_Kernel.vhd:1172:93  */
  assign n1365_o = n1364_o & n1362_o;
  /* TG68KdotC_Kernel.vhd:1172:127  */
  assign n1367_o = set_rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1172:113  */
  assign n1368_o = n1365_o | n1367_o;
  /* TG68KdotC_Kernel.vhd:1172:164  */
  assign n1369_o = ~interrupt;
  /* TG68KdotC_Kernel.vhd:1172:151  */
  assign n1370_o = n1369_o & stop;
  /* TG68KdotC_Kernel.vhd:1172:138  */
  assign n1371_o = n1368_o | n1370_o;
  /* TG68KdotC_Kernel.vhd:1172:181  */
  assign n1372_o = set_exec[31];
  /* TG68KdotC_Kernel.vhd:1172:170  */
  assign n1373_o = n1371_o | n1372_o;
  /* TG68KdotC_Kernel.vhd:1176:59  */
  assign n1374_o = exec_write_back & execopc;
  /* TG68KdotC_Kernel.vhd:1184:60  */
  assign n1377_o = setstate == 2'b01;
  /* TG68KdotC_Kernel.vhd:1187:59  */
  assign n1378_o = exec[29];
  /* TG68KdotC_Kernel.vhd:1191:58  */
  assign n1379_o = set[73];
  /* TG68KdotC_Kernel.vhd:1196:67  */
  assign n1381_o = set_datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:1196:85  */
  assign n1382_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1196:73  */
  assign n1383_o = n1382_o & n1381_o;
  /* TG68KdotC_Kernel.vhd:1199:63  */
  assign n1384_o = set[72];
  /* TG68KdotC_Kernel.vhd:1199:57  */
  assign n1387_o = n1384_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1196:49  */
  assign n1390_o = n1383_o ? 6'b101111 : 6'b100111;
  /* TG68KdotC_Kernel.vhd:1196:49  */
  assign n1393_o = n1383_o ? 6'b101111 : 6'b100111;
  /* TG68KdotC_Kernel.vhd:1196:49  */
  assign n1395_o = n1383_o ? n1387_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1191:49  */
  assign n1397_o = n1379_o ? 6'b100001 : n1390_o;
  /* TG68KdotC_Kernel.vhd:1191:49  */
  assign n1399_o = n1379_o ? 6'b100001 : n1393_o;
  /* TG68KdotC_Kernel.vhd:1191:49  */
  assign n1401_o = n1379_o ? 1'b0 : n1395_o;
  /* TG68KdotC_Kernel.vhd:1187:49  */
  assign n1402_o = n1378_o ? set_memmask : n1397_o;
  /* TG68KdotC_Kernel.vhd:1187:49  */
  assign n1403_o = n1378_o ? set_memmask : n1399_o;
  /* TG68KdotC_Kernel.vhd:1187:49  */
  assign n1404_o = n1378_o ? set_oddout : n1401_o;
  /* TG68KdotC_Kernel.vhd:1184:49  */
  assign n1406_o = n1377_o ? 6'b111111 : n1402_o;
  /* TG68KdotC_Kernel.vhd:1184:49  */
  assign n1408_o = n1377_o ? 6'b111111 : n1403_o;
  /* TG68KdotC_Kernel.vhd:1184:49  */
  assign n1409_o = n1377_o ? oddout : n1404_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1410_o = n1374_o ? 2'b01 : n1346_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1412_o = n1374_o ? 2'b11 : setstate;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1414_o = n1374_o ? 1'b0 : setaddrvalue;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1415_o = n1374_o ? wbmemmask : n1406_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1416_o = n1374_o ? wbmemmask : n1408_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1417_o = n1374_o ? oddout : n1409_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1418_o = n1373_o ? n1346_o : n1410_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1420_o = n1373_o ? 2'b01 : n1412_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1422_o = n1373_o ? 1'b0 : n1414_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1424_o = n1373_o ? 6'b111111 : n1415_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1425_o = n1373_o ? wbmemmask : n1416_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1426_o = n1373_o ? oddout : n1417_o;
  /* TG68KdotC_Kernel.vhd:1215:78  */
  assign n1427_o = set_writepcbig | writepcbig;
  /* TG68KdotC_Kernel.vhd:1211:41  */
  assign n1429_o = decodeopc ? 1'b0 : n1427_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1430_o = n1488_o ? set_rot_bits : rot_bits;
  /* TG68KdotC_Kernel.vhd:1217:65  */
  assign n1431_o = exec[24];
  /* TG68KdotC_Kernel.vhd:1217:58  */
  assign n1432_o = decodeopc | n1431_o;
  /* TG68KdotC_Kernel.vhd:1217:92  */
  assign n1434_o = rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1217:82  */
  assign n1435_o = n1432_o | n1434_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1436_o = n1489_o ? set_rot_cnt : rot_cnt;
  /* TG68KdotC_Kernel.vhd:1223:55  */
  assign n1437_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1223:86  */
  assign n1438_o = set[62];
  /* TG68KdotC_Kernel.vhd:1223:79  */
  assign n1439_o = n1438_o & ea_only;
  /* TG68KdotC_Kernel.vhd:1223:63  */
  assign n1440_o = n1437_o | n1439_o;
  /* TG68KdotC_Kernel.vhd:1223:41  */
  assign n1442_o = n1440_o ? 1'b0 : suppress_base;
  /* TG68KdotC_Kernel.vhd:1221:41  */
  assign n1444_o = set_suppress_base ? 1'b1 : n1442_o;
  /* TG68KdotC_Kernel.vhd:1227:57  */
  assign n1445_o = state[1];
  /* TG68KdotC_Kernel.vhd:1230:75  */
  assign n1446_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:1227:49  */
  assign n1447_o = n1445_o ? last_opc_read : n1446_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1448_o = n1482_o ? n1447_o : brief;
  /* TG68KdotC_Kernel.vhd:1234:66  */
  assign n1449_o = ~berr;
  /* TG68KdotC_Kernel.vhd:1234:58  */
  assign n1450_o = n1449_o & setopcode;
  /* TG68KdotC_Kernel.vhd:1235:57  */
  assign n1452_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1236:76  */
  assign n1453_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:1235:49  */
  assign n1454_o = n1452_o ? n1453_o : last_opc_read;
  /* TG68KdotC_Kernel.vhd:1235:49  */
  assign n1455_o = n1452_o ? tg68_pc : last_opc_pc;
  /* TG68KdotC_Kernel.vhd:1243:64  */
  assign n1456_o = setinterrupt | setopcode;
  /* TG68KdotC_Kernel.vhd:1248:68  */
  assign n1457_o = setnextpass | regdirectsource;
  /* TG68KdotC_Kernel.vhd:1248:49  */
  assign n1459_o = n1457_o ? 1'b1 : nextpass;
  /* TG68KdotC_Kernel.vhd:1243:41  */
  assign n1461_o = n1456_o ? 16'b0100111001110001 : opcode;
  /* TG68KdotC_Kernel.vhd:1243:41  */
  assign n1463_o = n1456_o ? 1'b0 : n1459_o;
  /* TG68KdotC_Kernel.vhd:1234:41  */
  assign n1464_o = n1450_o ? n1454_o : n1461_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1465_o = n1477_o ? n1455_o : exe_pc;
  /* TG68KdotC_Kernel.vhd:1234:41  */
  assign n1467_o = n1450_o ? 1'b0 : n1463_o;
  /* TG68KdotC_Kernel.vhd:1253:58  */
  assign n1468_o = decodeopc | interrupt;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1469_o = n1493_o ? flagssr : trap_sr;
  assign n1470_o = n9925_o[1:0];
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1471_o = clkena_lw ? n1418_o : n1470_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1472_o = clkena_lw ? n1420_o : state;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1473_o = clkena_lw ? set_datatype : exe_datatype;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1474_o = clkena_lw ? n1422_o : addrvalue;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1475_o = clkena_lw ? n1464_o : opcode;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1476_o = clkena_lw ? opcode : exe_opcode;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1477_o = n1450_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1478_o = n1302_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1479_o = n1302_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1480_o = clkena_lw ? n1467_o : nextpass;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1481_o = clkena_lw ? n1317_o : tg68_pc_word;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1482_o = getbrief & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1483_o = clkena_lw ? n1357_o : exec_write_back;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1484_o = clkena_lw ? n1429_o : writepcbig;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1485_o = clkena_lw ? setopcode : decodeopc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1486_o = clkena_lw ? setexecopc : execopc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1487_o = clkena_lw ? setendopc : endopc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1488_o = decodeopc & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1489_o = n1435_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1490_o = clkena_lw ? n1319_o : trap_berr;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1491_o = clkena_lw ? n1321_o : trap_trace;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1492_o = clkena_lw ? n1323_o : trap_interrupt;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1493_o = n1468_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1494_o = clkena_lw ? n1292_o : make_berr;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1495_o = clkena_lw ? n1265_o : stop;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1496_o = setinterrupt & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1497_o = clkena_lw ? n1300_o : ipl_vec;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1498_o = clkena_lw ? setinterrupt : interrupt;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1499_o = clkena_lw ? n1444_o : suppress_base;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1500_o = clkena_lw ? n1424_o : n1257_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1502_o = clkena_lw ? 4'b1111 : n1258_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1503_o = clkena_lw ? n1425_o : wbmemmask;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1504_o = clkena_lw ? n1426_o : oddout;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1505_o = n1324_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1506_o = n1324_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1507_o = n1324_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1508_o = n1324_o & clkena_lw;
  assign n1509_o = n9925_o[1:0];
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1510_o = reset ? n1509_o : n1471_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1512_o = reset ? 32'b00000000000000000000000000000100 : n1256_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1514_o = reset ? 2'b01 : n1472_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1515_o = reset ? exe_datatype : n1473_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1517_o = reset ? 1'b0 : n1474_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1519_o = reset ? 16'b0010111001111001 : n1475_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1520_o = reset ? exe_opcode : n1476_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1521_o = reset ? exe_pc : n1465_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1522_o = reset ? last_opc_pc : n1304_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1524_o = reset ? 16'b0100111011111001 : n1305_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1525_o = reset ? nextpass : n1480_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1527_o = reset ? 1'b0 : n1481_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1528_o = reset ? brief : n1448_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1530_o = reset ? 1'b0 : n1483_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1532_o = reset ? 1'b0 : n1484_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1534_o = reset ? 1'b0 : n1485_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1536_o = reset ? 1'b0 : n1486_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1538_o = reset ? 1'b0 : n1487_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1539_o = reset ? rot_bits : n1430_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1541_o = reset ? 6'b000001 : n1436_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1543_o = reset ? 1'b0 : n1490_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1545_o = reset ? 1'b0 : n1491_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1547_o = reset ? 1'b0 : n1492_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1548_o = reset ? trap_sr : n1469_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1550_o = reset ? 1'b0 : n1494_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1552_o = reset ? 1'b0 : n1495_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1553_o = reset ? ripl_nr : n1293_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1554_o = reset ? ipl_vec : n1497_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1556_o = reset ? 1'b0 : n1498_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1558_o = reset ? 1'b0 : n1499_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1560_o = reset ? 6'b111111 : n1500_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1561_o = reset ? memread : n1502_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1562_o = reset ? wbmemmask : n1503_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1563_o = reset ? oddout : n1504_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1564_o = reset ? alu_width : n1329_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1565_o = reset ? alu_bf_shift : n1330_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1566_o = reset ? alu_bf_ffo_offset : n1331_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1567_o = reset ? alu_bf_loffset : n1332_o;
  /* TG68KdotC_Kernel.vhd:1264:54  */
  assign n1608_o = set_pcbase | pcbase;
  /* TG68KdotC_Kernel.vhd:1265:60  */
  assign n1609_o = state[1];
  /* TG68KdotC_Kernel.vhd:1265:81  */
  assign n1610_o = ~movem_run;
  /* TG68KdotC_Kernel.vhd:1265:68  */
  assign n1611_o = n1610_o & n1609_o;
  /* TG68KdotC_Kernel.vhd:1265:51  */
  assign n1612_o = setexecopc | n1611_o;
  /* TG68KdotC_Kernel.vhd:1265:33  */
  assign n1614_o = n1612_o ? 1'b0 : n1608_o;
  /* TG68KdotC_Kernel.vhd:1263:25  */
  assign n1615_o = clkena_lw ? n1614_o : pcbase;
  /* TG68KdotC_Kernel.vhd:1261:25  */
  assign n1617_o = reset ? 1'b1 : n1615_o;
  /* TG68KdotC_Kernel.vhd:1271:54  */
  assign n1618_o = set[0];
  /* TG68KdotC_Kernel.vhd:1271:70  */
  assign n1619_o = set[85];
  /* TG68KdotC_Kernel.vhd:1271:64  */
  assign n1620_o = n1618_o | n1619_o;
  /* TG68KdotC_Kernel.vhd:1272:58  */
  assign n1623_o = set[3];
  /* TG68KdotC_Kernel.vhd:1272:73  */
  assign n1624_o = set[86];
  /* TG68KdotC_Kernel.vhd:1272:67  */
  assign n1625_o = n1623_o | n1624_o;
  assign n1626_o = set[88:87];
  /* TG68KdotC_Kernel.vhd:1274:52  */
  assign n1627_o = set[47];
  /* TG68KdotC_Kernel.vhd:1274:67  */
  assign n1628_o = set[48];
  /* TG68KdotC_Kernel.vhd:1274:61  */
  assign n1629_o = n1627_o | n1628_o;
  assign n1630_o = set[84:49];
  assign n1631_o = set[47:0];
  /* TG68KdotC_Kernel.vhd:1276:58  */
  assign n1632_o = set_exec | set;
  /* TG68KdotC_Kernel.vhd:1277:67  */
  assign n1633_o = set_exec[0];
  /* TG68KdotC_Kernel.vhd:1277:83  */
  assign n1634_o = set[0];
  /* TG68KdotC_Kernel.vhd:1277:77  */
  assign n1635_o = n1633_o | n1634_o;
  /* TG68KdotC_Kernel.vhd:1277:99  */
  assign n1636_o = set[85];
  /* TG68KdotC_Kernel.vhd:1277:93  */
  assign n1637_o = n1635_o | n1636_o;
  assign n1639_o = n1632_o[84:0];
  /* TG68KdotC_Kernel.vhd:1278:71  */
  assign n1640_o = set_exec[3];
  /* TG68KdotC_Kernel.vhd:1278:86  */
  assign n1641_o = set[3];
  /* TG68KdotC_Kernel.vhd:1278:80  */
  assign n1642_o = n1640_o | n1641_o;
  /* TG68KdotC_Kernel.vhd:1278:101  */
  assign n1643_o = set[86];
  /* TG68KdotC_Kernel.vhd:1278:95  */
  assign n1644_o = n1642_o | n1643_o;
  assign n1645_o = n1632_o[88:87];
  /* TG68KdotC_Kernel.vhd:1275:33  */
  assign n1647_o = setexecopc ? set_exec_tas : 1'b0;
  assign n1649_o = {n1645_o, n1644_o, n1637_o, n1639_o};
  assign n1650_o = {n1626_o, n1625_o, n1620_o, n1630_o, n1629_o, n1631_o};
  /* TG68KdotC_Kernel.vhd:1281:56  */
  assign n1652_o = set[71];
  /* TG68KdotC_Kernel.vhd:1281:69  */
  assign n1653_o = n1652_o | setopcode;
  assign n1654_o = n1649_o[88:72];
  assign n1655_o = n1650_o[88:72];
  /* TG68KdotC_Kernel.vhd:1275:33  */
  assign n1656_o = setexecopc ? n1654_o : n1655_o;
  assign n1657_o = n1649_o[70:0];
  assign n1658_o = n1650_o[70:0];
  /* TG68KdotC_Kernel.vhd:1275:33  */
  assign n1659_o = setexecopc ? n1657_o : n1658_o;
  assign n1661_o = {n1656_o, n1653_o, n1659_o};
  /* TG68KdotC_Kernel.vhd:1291:26  */
  assign n1669_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:1292:48  */
  assign n1670_o = reg_qa[4:0];
  /* TG68KdotC_Kernel.vhd:1292:41  */
  assign n1672_o = {1'b0, n1670_o};
  /* TG68KdotC_Kernel.vhd:1294:48  */
  assign n1673_o = sndopc[10:6];
  /* TG68KdotC_Kernel.vhd:1294:41  */
  assign n1675_o = {1'b0, n1673_o};
  /* TG68KdotC_Kernel.vhd:1296:26  */
  assign n1677_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:1300:61  */
  assign n1678_o = sndopc[10:6];
  assign n1680_o = n1679_o[31:5];
  assign n1681_o = {n1680_o, n1678_o};
  /* TG68KdotC_Kernel.vhd:1296:17  */
  assign n1682_o = n1677_o ? reg_qa : n1681_o;
  /* TG68KdotC_Kernel.vhd:1304:26  */
  assign n1684_o = sndopc[5];
  /* TG68KdotC_Kernel.vhd:1305:55  */
  assign n1685_o = reg_qb[4:0];
  /* TG68KdotC_Kernel.vhd:1305:67  */
  assign n1687_o = n1685_o - 5'b00001;
  /* TG68KdotC_Kernel.vhd:1307:55  */
  assign n1688_o = sndopc[4:0];
  /* TG68KdotC_Kernel.vhd:1307:67  */
  assign n1690_o = n1688_o - 5'b00001;
  /* TG68KdotC_Kernel.vhd:1304:17  */
  assign n1691_o = n1684_o ? n1687_o : n1690_o;
  /* TG68KdotC_Kernel.vhd:1309:37  */
  assign n1692_o = bf_width + bf_offset;
  /* TG68KdotC_Kernel.vhd:1310:43  */
  assign n1693_o = bf_bhits[3];
  /* TG68KdotC_Kernel.vhd:1310:31  */
  assign n1694_o = ~n1693_o;
  /* TG68KdotC_Kernel.vhd:1314:26  */
  assign n1695_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:1314:39  */
  assign n1697_o = n1695_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1315:41  */
  assign n1699_o = 6'b100000 - bf_shift;
  assign n1702_o = n1699_o[4:0];
  assign n1703_o = bf_shift[4:0];
  /* TG68KdotC_Kernel.vhd:1314:17  */
  assign n1704_o = n1697_o ? n1702_o : n1703_o;
  /* TG68KdotC_Kernel.vhd:1321:26  */
  assign n1705_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:1321:38  */
  assign n1707_o = n1705_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1322:34  */
  assign n1708_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:1322:47  */
  assign n1710_o = n1708_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1323:53  */
  assign n1712_o = bf_bhits + 6'b000001;
  /* TG68KdotC_Kernel.vhd:1325:47  */
  assign n1714_o = 6'b011111 - bf_bhits;
  assign n1717_o = n1712_o[4:0];
  assign n1718_o = n1714_o[4:0];
  /* TG68KdotC_Kernel.vhd:1322:25  */
  assign n1719_o = n1710_o ? n1717_o : n1718_o;
  /* TG68KdotC_Kernel.vhd:1329:34  */
  assign n1720_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:1329:47  */
  assign n1722_o = n1720_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1330:69  */
  assign n1723_o = bf_bhits[2:0];
  /* TG68KdotC_Kernel.vhd:1330:60  */
  assign n1725_o = {3'b000, n1723_o};
  /* TG68KdotC_Kernel.vhd:1330:53  */
  assign n1727_o = 6'b011001 + n1725_o;
  assign n1729_o = n1727_o[4:0];
  /* TG68KdotC_Kernel.vhd:1333:66  */
  assign n1730_o = bf_bhits[2:0];
  /* TG68KdotC_Kernel.vhd:1333:57  */
  assign n1732_o = 3'b111 - n1730_o;
  /* TG68KdotC_Kernel.vhd:1333:50  */
  assign n1734_o = {3'b000, n1732_o};
  assign n1735_o = {1'b0, n1729_o};
  /* TG68KdotC_Kernel.vhd:1329:25  */
  assign n1736_o = n1722_o ? n1735_o : n1734_o;
  assign n1738_o = n1672_o[4:3];
  assign n1739_o = n1675_o[4:3];
  /* TG68KdotC_Kernel.vhd:1291:17  */
  assign n1740_o = n1669_o ? n1738_o : n1739_o;
  /* TG68KdotC_Kernel.vhd:1321:17  */
  assign n1741_o = n1707_o ? n1740_o : 2'b00;
  assign n1742_o = n1672_o[5];
  assign n1743_o = n1675_o[5];
  /* TG68KdotC_Kernel.vhd:1291:17  */
  assign n1744_o = n1669_o ? n1742_o : n1743_o;
  assign n1745_o = n1672_o[2:0];
  assign n1746_o = n1675_o[2:0];
  /* TG68KdotC_Kernel.vhd:1291:17  */
  assign n1747_o = n1669_o ? n1745_o : n1746_o;
  assign n1748_o = {1'b0, n1719_o};
  /* TG68KdotC_Kernel.vhd:1321:17  */
  assign n1749_o = n1707_o ? n1748_o : n1736_o;
  /* TG68KdotC_Kernel.vhd:1338:30  */
  assign n1750_o = bf_bhits[5:3];
  /* TG68KdotC_Kernel.vhd:1339:25  */
  assign n1752_o = n1750_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1341:25  */
  assign n1754_o = n1750_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1343:25  */
  assign n1756_o = n1750_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1345:25  */
  assign n1758_o = n1750_o == 3'b011;
  assign n1759_o = {n1758_o, n1756_o, n1754_o, n1752_o};
  /* TG68KdotC_Kernel.vhd:1338:17  */
  always @*
    case (n1759_o)
      4'b1000: n1765_o = 6'b100001;
      4'b0100: n1765_o = 6'b100011;
      4'b0010: n1765_o = 6'b100111;
      4'b0001: n1765_o = 6'b101111;
      default: n1765_o = 6'b100000;
    endcase
  /* TG68KdotC_Kernel.vhd:1350:28  */
  assign n1767_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1350:17  */
  assign n1769_o = n1767_o ? 6'b100111 : n1765_o;
  /* TG68KdotC_Kernel.vhd:1360:24  */
  assign n1773_o = exec[17];
  /* TG68KdotC_Kernel.vhd:1361:59  */
  assign n1774_o = last_data_read[15:8];
  /* TG68KdotC_Kernel.vhd:1361:41  */
  assign n1775_o = flagssr & n1774_o;
  /* TG68KdotC_Kernel.vhd:1362:27  */
  assign n1776_o = exec[18];
  /* TG68KdotC_Kernel.vhd:1363:59  */
  assign n1777_o = last_data_read[15:8];
  /* TG68KdotC_Kernel.vhd:1363:41  */
  assign n1778_o = flagssr ^ n1777_o;
  /* TG68KdotC_Kernel.vhd:1364:27  */
  assign n1779_o = exec[19];
  /* TG68KdotC_Kernel.vhd:1365:58  */
  assign n1780_o = last_data_read[15:8];
  /* TG68KdotC_Kernel.vhd:1365:41  */
  assign n1781_o = flagssr | n1780_o;
  /* TG68KdotC_Kernel.vhd:1367:39  */
  assign n1782_o = op2out[15:8];
  /* TG68KdotC_Kernel.vhd:1364:17  */
  assign n1783_o = n1779_o ? n1781_o : n1782_o;
  /* TG68KdotC_Kernel.vhd:1362:17  */
  assign n1784_o = n1776_o ? n1778_o : n1783_o;
  /* TG68KdotC_Kernel.vhd:1360:17  */
  assign n1785_o = n1773_o ? n1775_o : n1784_o;
  /* TG68KdotC_Kernel.vhd:1379:62  */
  assign n1788_o = flagssr[7];
  /* TG68KdotC_Kernel.vhd:1380:47  */
  assign n1789_o = set[41];
  /* TG68KdotC_Kernel.vhd:1381:59  */
  assign n1790_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:1380:41  */
  assign n1791_o = n1789_o ? n1790_o : presvmode;
  /* TG68KdotC_Kernel.vhd:1378:33  */
  assign n1792_o = setopcode ? n1788_o : make_trace;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1793_o = n1880_o ? n1791_o : svmode;
  /* TG68KdotC_Kernel.vhd:1386:50  */
  assign n1794_o = trap_berr | trap_illegal;
  /* TG68KdotC_Kernel.vhd:1386:70  */
  assign n1795_o = n1794_o | trap_addr_error;
  /* TG68KdotC_Kernel.vhd:1386:93  */
  assign n1796_o = n1795_o | trap_priv;
  /* TG68KdotC_Kernel.vhd:1386:110  */
  assign n1797_o = n1796_o | trap_1010;
  /* TG68KdotC_Kernel.vhd:1386:127  */
  assign n1798_o = n1797_o | trap_1111;
  assign n1800_o = flagssr[7];
  /* TG68KdotC_Kernel.vhd:1386:33  */
  assign n1801_o = n1798_o ? 1'b0 : n1800_o;
  /* TG68KdotC_Kernel.vhd:1386:33  */
  assign n1803_o = n1798_o ? 1'b0 : n1792_o;
  /* TG68KdotC_Kernel.vhd:1390:39  */
  assign n1804_o = set[41];
  /* TG68KdotC_Kernel.vhd:1391:54  */
  assign n1805_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1392:55  */
  assign n1806_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1393:50  */
  assign n1807_o = ~presvmode;
  assign n1808_o = n9925_o[2];
  /* TG68KdotC_Kernel.vhd:1390:33  */
  assign n1809_o = n1804_o ? n1807_o : n1808_o;
  assign n1810_o = flagssr[5];
  /* TG68KdotC_Kernel.vhd:1390:33  */
  assign n1811_o = n1804_o ? n1806_o : n1810_o;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1812_o = n1881_o ? n1805_o : presvmode;
  /* TG68KdotC_Kernel.vhd:1395:47  */
  assign n1814_o = micro_state == 7'b0110110;
  /* TG68KdotC_Kernel.vhd:1395:33  */
  assign n1816_o = n1814_o ? 1'b0 : n1801_o;
  /* TG68KdotC_Kernel.vhd:1398:60  */
  assign n1818_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1398:51  */
  assign n1819_o = n1818_o & trap_trace;
  /* TG68KdotC_Kernel.vhd:1398:33  */
  assign n1821_o = n1819_o ? 1'b0 : n1803_o;
  /* TG68KdotC_Kernel.vhd:1401:40  */
  assign n1822_o = exec[59];
  /* TG68KdotC_Kernel.vhd:1401:55  */
  assign n1823_o = n1822_o | set_stop;
  assign n1825_o = flagssr[4:0];
  assign n1826_o = flagssr[6];
  assign n1827_o = {n1816_o, n1826_o, n1811_o, n1825_o};
  /* TG68KdotC_Kernel.vhd:1404:50  */
  assign n1829_o = trap_interrupt & interrupt;
  assign n1830_o = data_read[10:8];
  assign n1831_o = n1827_o[2:0];
  /* TG68KdotC_Kernel.vhd:1401:33  */
  assign n1832_o = n1823_o ? n1830_o : n1831_o;
  /* TG68KdotC_Kernel.vhd:1404:33  */
  assign n1833_o = n1829_o ? ripl_nr : n1832_o;
  assign n1834_o = data_read[15:11];
  assign n1835_o = n1827_o[7:3];
  /* TG68KdotC_Kernel.vhd:1401:33  */
  assign n1836_o = n1823_o ? n1834_o : n1835_o;
  /* TG68KdotC_Kernel.vhd:1407:40  */
  assign n1837_o = exec[52];
  /* TG68KdotC_Kernel.vhd:1409:54  */
  assign n1838_o = srin[5];
  /* TG68KdotC_Kernel.vhd:1410:43  */
  assign n1839_o = exec[35];
  /* TG68KdotC_Kernel.vhd:1411:57  */
  assign n1840_o = flagssr[5];
  /* TG68KdotC_Kernel.vhd:1410:33  */
  assign n1841_o = n1839_o ? n1840_o : n1809_o;
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1842_o = n1837_o ? n1838_o : n1841_o;
  assign n1843_o = {n1836_o, n1833_o};
  /* TG68KdotC_Kernel.vhd:1413:33  */
  assign n1846_o = interrupt ? 1'b1 : n1842_o;
  /* TG68KdotC_Kernel.vhd:1416:39  */
  assign n1847_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1416:42  */
  assign n1848_o = ~n1847_o;
  assign n1851_o = srin[4];
  assign n1852_o = n1843_o[4];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1853_o = n1837_o ? n1851_o : n1852_o;
  /* TG68KdotC_Kernel.vhd:1416:33  */
  assign n1854_o = n1848_o ? 1'b0 : n1853_o;
  assign n1855_o = srin[6];
  assign n1856_o = n1843_o[6];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1857_o = n1837_o ? n1855_o : n1856_o;
  /* TG68KdotC_Kernel.vhd:1416:33  */
  assign n1858_o = n1848_o ? 1'b0 : n1857_o;
  assign n1865_o = srin[7];
  assign n1866_o = n1843_o[7];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1867_o = n1837_o ? n1865_o : n1866_o;
  assign n1868_o = srin[5];
  assign n1869_o = n1843_o[5];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1870_o = n1837_o ? n1868_o : n1869_o;
  assign n1872_o = srin[2:0];
  assign n1873_o = n1843_o[2:0];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1874_o = n1837_o ? n1872_o : n1873_o;
  assign n1875_o = n9925_o[2];
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1876_o = clkena_lw ? n1846_o : n1875_o;
  assign n1877_o = {n1867_o, n1858_o, n1870_o, n1854_o, 1'b0, n1874_o};
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1878_o = clkena_lw ? n1877_o : flagssr;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1879_o = clkena_lw ? n1821_o : make_trace;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1880_o = setopcode & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1881_o = n1804_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1882_o = reset ? 1'b1 : n1876_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1884_o = reset ? 8'b00100111 : n1878_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1886_o = reset ? 1'b0 : n1879_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1888_o = reset ? 1'b1 : n1793_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1890_o = reset ? 1'b1 : n1812_o;
  /* TG68KdotC_Kernel.vhd:1453:39  */
  assign n1900_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:1495:27  */
  assign n1902_o = rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1496:47  */
  assign n1904_o = rot_cnt - 6'b000001;
  /* TG68KdotC_Kernel.vhd:1495:17  */
  assign n1906_o = n1902_o ? n1904_o : 6'b000001;
  /* TG68KdotC_Kernel.vhd:1507:28  */
  assign n1912_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1508:25  */
  assign n1914_o = n1912_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1509:25  */
  assign n1916_o = n1912_o == 2'b01;
  assign n1917_o = {n1916_o, n1914_o};
  /* TG68KdotC_Kernel.vhd:1507:17  */
  always @*
    case (n1917_o)
      2'b10: n1921_o = 2'b01;
      2'b01: n1921_o = 2'b00;
      default: n1921_o = 2'b10;
    endcase
  /* TG68KdotC_Kernel.vhd:1513:32  */
  assign n1922_o = exec_write_back & execopc;
  assign n1924_o = n1909_o[83];
  /* TG68KdotC_Kernel.vhd:1513:17  */
  assign n1925_o = n1922_o ? 1'b1 : n1924_o;
  /* TG68KdotC_Kernel.vhd:1517:34  */
  assign n1928_o = trap_berr & interrupt;
  /* TG68KdotC_Kernel.vhd:1519:37  */
  assign n1929_o = ~presvmode;
  assign n1931_o = n1909_o[41];
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1932_o = n1938_o ? 1'b1 : n1931_o;
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1935_o = n1928_o ? 2'b01 : 2'b00;
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1938_o = n1929_o & n1928_o;
  assign n1940_o = n1909_o[40:39];
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1943_o = n1928_o ? 7'b1000110 : 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1524:42  */
  assign n1945_o = ~trapd;
  /* TG68KdotC_Kernel.vhd:1524:33  */
  assign n1946_o = n1945_o & trapmake;
  /* TG68KdotC_Kernel.vhd:1525:31  */
  assign n1947_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1525:59  */
  assign n1948_o = trap_trapv | set_z_error;
  /* TG68KdotC_Kernel.vhd:1525:85  */
  assign n1949_o = exec[43];
  /* TG68KdotC_Kernel.vhd:1525:78  */
  assign n1950_o = n1948_o | n1949_o;
  /* TG68KdotC_Kernel.vhd:1525:39  */
  assign n1951_o = n1950_o & n1947_o;
  /* TG68KdotC_Kernel.vhd:1527:25  */
  assign n1954_o = trap_addr_error ? 7'b1000110 : 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1525:25  */
  assign n1956_o = n1951_o ? 7'b0110010 : n1954_o;
  /* TG68KdotC_Kernel.vhd:1532:46  */
  assign n1957_o = ~use_vbr_stackframe;
  assign n1959_o = n1909_o[25];
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1960_o = n1967_o ? 1'b1 : n1959_o;
  /* TG68KdotC_Kernel.vhd:1536:37  */
  assign n1961_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1963_o = n1968_o ? 1'b1 : n1932_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1965_o = n1946_o ? 2'b01 : n1935_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1967_o = n1957_o & n1946_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1968_o = n1961_o & n1946_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1971_o = n1946_o ? n1956_o : n1943_o;
  /* TG68KdotC_Kernel.vhd:1541:31  */
  assign n1973_o = micro_state == 7'b0100111;
  /* TG68KdotC_Kernel.vhd:1541:55  */
  assign n1974_o = trap_trace & interrupt;
  /* TG68KdotC_Kernel.vhd:1541:37  */
  assign n1975_o = n1973_o | n1974_o;
  /* TG68KdotC_Kernel.vhd:1543:50  */
  assign n1976_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1543:43  */
  assign n1977_o = n1976_o & trap_trace;
  /* TG68KdotC_Kernel.vhd:1543:25  */
  assign n1980_o = n1977_o ? 7'b0110010 : 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1553:37  */
  assign n1981_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1983_o = n1986_o ? 1'b1 : n1963_o;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1985_o = n1975_o ? 2'b01 : n1965_o;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1986_o = n1981_o & n1975_o;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1987_o = n1975_o ? n1980_o : n1971_o;
  /* TG68KdotC_Kernel.vhd:1558:24  */
  assign n1989_o = micro_state == 7'b0100111;
  /* TG68KdotC_Kernel.vhd:1558:51  */
  assign n1990_o = trap_trace & interrupt;
  /* TG68KdotC_Kernel.vhd:1558:31  */
  assign n1991_o = n1989_o | n1990_o;
  /* TG68KdotC_Kernel.vhd:1559:24  */
  assign n1992_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1558:9  */
  assign n1994_o = n1997_o ? 1'b1 : n1983_o;
  /* TG68KdotC_Kernel.vhd:1558:9  */
  assign n1996_o = n1991_o ? 2'b01 : n1985_o;
  /* TG68KdotC_Kernel.vhd:1558:9  */
  assign n1997_o = n1992_o & n1991_o;
  /* TG68KdotC_Kernel.vhd:1565:46  */
  assign n1998_o = flagssr[5];
  /* TG68KdotC_Kernel.vhd:1565:49  */
  assign n1999_o = n1998_o != presvmode;
  /* TG68KdotC_Kernel.vhd:1565:35  */
  assign n2000_o = n1999_o & setexecopc;
  /* TG68KdotC_Kernel.vhd:1565:17  */
  assign n2002_o = n2000_o ? 1'b1 : n1994_o;
  /* TG68KdotC_Kernel.vhd:1571:34  */
  assign n2003_o = trap_interrupt & interrupt;
  /* TG68KdotC_Kernel.vhd:1571:17  */
  assign n2006_o = n2003_o ? 2'b10 : n1996_o;
  /* TG68KdotC_Kernel.vhd:1571:17  */
  assign n2007_o = n2003_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1571:17  */
  assign n2009_o = n2003_o ? 7'b0100111 : n1987_o;
  /* TG68KdotC_Kernel.vhd:1578:23  */
  assign n2010_o = set[41];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n2015_o = n2010_o ? 1'b1 : 1'b0;
  assign n2017_o = {1'b1, 1'b1};
  assign n2018_o = n1909_o[66:65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n2019_o = n2010_o ? n2017_o : n2018_o;
  /* TG68KdotC_Kernel.vhd:1584:27  */
  assign n2022_o = ~ea_only;
  /* TG68KdotC_Kernel.vhd:1584:39  */
  assign n2023_o = set[62];
  /* TG68KdotC_Kernel.vhd:1584:32  */
  assign n2024_o = n2023_o & n2022_o;
  /* TG68KdotC_Kernel.vhd:1584:17  */
  assign n2026_o = n2024_o ? 2'b10 : n2006_o;
  /* TG68KdotC_Kernel.vhd:1590:28  */
  assign n2027_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1590:52  */
  assign n2028_o = set_datatype[1];
  /* TG68KdotC_Kernel.vhd:1590:36  */
  assign n2029_o = n2028_o & n2027_o;
  assign n2031_o = n1909_o[73];
  /* TG68KdotC_Kernel.vhd:1590:17  */
  assign n2032_o = n2029_o ? 1'b1 : n2031_o;
  /* TG68KdotC_Kernel.vhd:1594:38  */
  assign n2035_o = decodeopc & ea_build_now;
  /* TG68KdotC_Kernel.vhd:1594:64  */
  assign n2036_o = exec[42];
  /* TG68KdotC_Kernel.vhd:1594:57  */
  assign n2037_o = n2035_o | n2036_o;
  /* TG68KdotC_Kernel.vhd:1595:36  */
  assign n2038_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1599:50  */
  assign n2040_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:1601:58  */
  assign n2042_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1601:70  */
  assign n2044_o = n2042_o == 3'b111;
  assign n2046_o = n1909_o[50];
  /* TG68KdotC_Kernel.vhd:1599:41  */
  assign n2047_o = n2051_o ? 1'b1 : n2046_o;
  assign n2048_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1599:41  */
  assign n2049_o = n2040_o ? 1'b1 : n2048_o;
  /* TG68KdotC_Kernel.vhd:1599:41  */
  assign n2051_o = n2044_o & n2040_o;
  /* TG68KdotC_Kernel.vhd:1605:50  */
  assign n2052_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:1607:58  */
  assign n2054_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1607:70  */
  assign n2056_o = n2054_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1605:41  */
  assign n2058_o = n2061_o ? 1'b1 : n2047_o;
  assign n2059_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1605:41  */
  assign n2060_o = n2052_o ? 1'b1 : n2059_o;
  /* TG68KdotC_Kernel.vhd:1605:41  */
  assign n2061_o = n2056_o & n2052_o;
  /* TG68KdotC_Kernel.vhd:1596:33  */
  assign n2063_o = n2038_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1596:43  */
  assign n2065_o = n2038_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1596:43  */
  assign n2066_o = n2063_o | n2065_o;
  /* TG68KdotC_Kernel.vhd:1596:49  */
  assign n2068_o = n2038_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1596:49  */
  assign n2069_o = n2066_o | n2068_o;
  /* TG68KdotC_Kernel.vhd:1611:33  */
  assign n2071_o = n2038_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:1613:33  */
  assign n2073_o = n2038_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:1617:52  */
  assign n2074_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1618:49  */
  assign n2076_o = n2074_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1620:49  */
  assign n2079_o = n2074_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1623:49  */
  assign n2082_o = n2074_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1628:49  */
  assign n2085_o = n2074_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1637:68  */
  assign n2087_o = datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:1637:57  */
  assign n2089_o = n2087_o ? 1'b1 : n2032_o;
  /* TG68KdotC_Kernel.vhd:1634:49  */
  assign n2091_o = n2074_o == 3'b100;
  assign n2092_o = {n2091_o, n2085_o, n2082_o, n2079_o, n2076_o};
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2095_o = 1'b1;
      5'b01000: n2095_o = 1'b0;
      5'b00100: n2095_o = 1'b0;
      5'b00010: n2095_o = 1'b0;
      5'b00001: n2095_o = 1'b0;
      default: n2095_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2098_o = 1'b0;
      5'b01000: n2098_o = 1'b1;
      5'b00100: n2098_o = 1'b0;
      5'b00010: n2098_o = 1'b0;
      5'b00001: n2098_o = 1'b0;
      default: n2098_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2101_o = 1'b1;
      5'b01000: n2101_o = 1'b0;
      5'b00100: n2101_o = 1'b0;
      5'b00010: n2101_o = 1'b0;
      5'b00001: n2101_o = 1'b0;
      default: n2101_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2105_o = 1'b0;
      5'b01000: n2105_o = 1'b1;
      5'b00100: n2105_o = 1'b1;
      5'b00010: n2105_o = 1'b0;
      5'b00001: n2105_o = 1'b0;
      default: n2105_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2109_o = 1'b0;
      5'b01000: n2109_o = 1'b1;
      5'b00100: n2109_o = 1'b1;
      5'b00010: n2109_o = 1'b0;
      5'b00001: n2109_o = 1'b0;
      default: n2109_o = 1'b0;
    endcase
  assign n2110_o = n1909_o[22];
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2111_o = n2110_o;
      5'b01000: n2111_o = 1'b1;
      5'b00100: n2111_o = 1'b1;
      5'b00010: n2111_o = n2110_o;
      5'b00001: n2111_o = n2110_o;
      default: n2111_o = n2110_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2112_o = n2089_o;
      5'b01000: n2112_o = n2032_o;
      5'b00100: n2112_o = n2032_o;
      5'b00010: n2112_o = 1'b1;
      5'b00001: n2112_o = n2032_o;
      default: n2112_o = n2032_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2117_o = n2009_o;
      5'b01000: n2117_o = 7'b0000101;
      5'b00100: n2117_o = 7'b0000100;
      5'b00010: n2117_o = 7'b0000010;
      5'b00001: n2117_o = 7'b0000010;
      default: n2117_o = n2009_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1616:33  */
  assign n2119_o = n2038_o == 3'b111;
  assign n2120_o = {n2119_o, n2073_o, n2071_o, n2069_o};
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2123_o = n2095_o;
      4'b0100: n2123_o = 1'b0;
      4'b0010: n2123_o = 1'b0;
      4'b0001: n2123_o = 1'b1;
      default: n2123_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2126_o = n2098_o;
      4'b0100: n2126_o = 1'b1;
      4'b0010: n2126_o = 1'b0;
      4'b0001: n2126_o = 1'b0;
      default: n2126_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2128_o = n2101_o;
      4'b0100: n2128_o = 1'b0;
      4'b0010: n2128_o = 1'b0;
      4'b0001: n2128_o = 1'b0;
      default: n2128_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2130_o = n2105_o;
      4'b0100: n2130_o = 1'b0;
      4'b0010: n2130_o = 1'b0;
      4'b0001: n2130_o = 1'b0;
      default: n2130_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2132_o = n2109_o;
      4'b0100: n2132_o = 1'b0;
      4'b0010: n2132_o = 1'b0;
      4'b0001: n2132_o = 1'b0;
      default: n2132_o = 1'b0;
    endcase
  assign n2133_o = n1909_o[22];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2134_o = n2111_o;
      4'b0100: n2134_o = n2133_o;
      4'b0010: n2134_o = n2133_o;
      4'b0001: n2134_o = n2133_o;
      default: n2134_o = n2133_o;
    endcase
  assign n2135_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2136_o = n2135_o;
      4'b0100: n2136_o = n2135_o;
      4'b0010: n2136_o = n2135_o;
      4'b0001: n2136_o = n2049_o;
      default: n2136_o = n2135_o;
    endcase
  assign n2137_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2138_o = n2137_o;
      4'b0100: n2138_o = n2137_o;
      4'b0010: n2138_o = n2137_o;
      4'b0001: n2138_o = n2060_o;
      default: n2138_o = n2137_o;
    endcase
  assign n2139_o = n1909_o[50];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2140_o = n2139_o;
      4'b0100: n2140_o = n2139_o;
      4'b0010: n2140_o = n2139_o;
      4'b0001: n2140_o = n2058_o;
      default: n2140_o = n2139_o;
    endcase
  assign n2141_o = n1909_o[62];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2142_o = n2141_o;
      4'b0100: n2142_o = n2141_o;
      4'b0010: n2142_o = n2141_o;
      4'b0001: n2142_o = 1'b1;
      default: n2142_o = n2141_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2143_o = n2112_o;
      4'b0100: n2143_o = n2032_o;
      4'b0010: n2143_o = n2032_o;
      4'b0001: n2143_o = n2032_o;
      default: n2143_o = n2032_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2146_o = n2117_o;
      4'b0100: n2146_o = 7'b0000101;
      4'b0010: n2146_o = 7'b0000100;
      4'b0001: n2146_o = n2009_o;
      default: n2146_o = n2009_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2148_o = n2037_o ? n2123_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2151_o = n2037_o ? n2126_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2154_o = n2037_o ? n2128_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2157_o = n2037_o ? n2130_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2160_o = n2037_o ? n2132_o : 1'b0;
  assign n2162_o = {n2138_o, n2136_o};
  assign n2163_o = n1909_o[22];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2164_o = n2037_o ? n2134_o : n2163_o;
  assign n2165_o = n1909_o[47:46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2166_o = n2037_o ? n2162_o : n2165_o;
  assign n2167_o = n1909_o[50];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2168_o = n2037_o ? n2140_o : n2167_o;
  assign n2169_o = n1909_o[62];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2170_o = n2037_o ? n2142_o : n2169_o;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2171_o = n2037_o ? n2143_o : n2032_o;
  assign n2177_o = n1909_o[49:48];
  assign n2178_o = n1909_o[64:63];
  assign n2179_o = n1909_o[61:51];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2180_o = n2037_o ? n2146_o : n2009_o;
  /* TG68KdotC_Kernel.vhd:1649:28  */
  assign n2181_o = tg68_pc[0];
  /* TG68KdotC_Kernel.vhd:1649:54  */
  assign n2183_o = micro_state == 7'b0000001;
  /* TG68KdotC_Kernel.vhd:1649:38  */
  assign n2184_o = n2183_o & n2181_o;
  /* TG68KdotC_Kernel.vhd:1653:28  */
  assign n2185_o = opcode[15:12];
  /* TG68KdotC_Kernel.vhd:1656:34  */
  assign n2186_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1656:52  */
  assign n2187_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1656:64  */
  assign n2189_o = n2187_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1656:42  */
  assign n2190_o = n2189_o & n2186_o;
  /* TG68KdotC_Kernel.vhd:1660:42  */
  assign n2193_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1660:45  */
  assign n2194_o = ~n2193_o;
  assign n2198_o = n1909_o[37];
  /* TG68KdotC_Kernel.vhd:1660:33  */
  assign n2199_o = n2194_o ? 1'b1 : n2198_o;
  /* TG68KdotC_Kernel.vhd:1660:33  */
  assign n2201_o = n2194_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1660:33  */
  assign n2203_o = n2194_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1666:50  */
  assign n2204_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2206_o = n2212_o ? 1'b1 : n2199_o;
  /* TG68KdotC_Kernel.vhd:1669:50  */
  assign n2207_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1669:53  */
  assign n2208_o = ~n2207_o;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2210_o = n2211_o ? 1'b1 : n2154_o;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2211_o = n2208_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2212_o = n2204_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2214_o = decodeopc ? 7'b1001010 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1674:33  */
  assign n2217_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1678:42  */
  assign n2218_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1678:59  */
  assign n2219_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1678:72  */
  assign n2221_o = n2219_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1678:50  */
  assign n2222_o = n2218_o | n2221_o;
  /* TG68KdotC_Kernel.vhd:1679:50  */
  assign n2223_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1679:62  */
  assign n2225_o = n2223_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1680:51  */
  assign n2226_o = opcode[8:3];
  /* TG68KdotC_Kernel.vhd:1680:63  */
  assign n2228_o = n2226_o != 6'b000111;
  /* TG68KdotC_Kernel.vhd:1680:83  */
  assign n2229_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:1680:86  */
  assign n2230_o = ~n2229_o;
  /* TG68KdotC_Kernel.vhd:1680:74  */
  assign n2231_o = n2228_o | n2230_o;
  /* TG68KdotC_Kernel.vhd:1679:70  */
  assign n2232_o = n2231_o & n2225_o;
  /* TG68KdotC_Kernel.vhd:1681:51  */
  assign n2233_o = opcode[8:2];
  /* TG68KdotC_Kernel.vhd:1681:63  */
  assign n2235_o = n2233_o != 7'b1001111;
  /* TG68KdotC_Kernel.vhd:1681:84  */
  assign n2236_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:1681:96  */
  assign n2238_o = n2236_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1681:75  */
  assign n2239_o = n2235_o | n2238_o;
  /* TG68KdotC_Kernel.vhd:1680:92  */
  assign n2240_o = n2239_o & n2232_o;
  /* TG68KdotC_Kernel.vhd:1682:51  */
  assign n2241_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1682:63  */
  assign n2243_o = n2241_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1682:78  */
  assign n2244_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1682:90  */
  assign n2246_o = n2244_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1682:69  */
  assign n2247_o = n2243_o | n2246_o;
  /* TG68KdotC_Kernel.vhd:1682:107  */
  assign n2248_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1682:119  */
  assign n2250_o = n2248_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1682:98  */
  assign n2251_o = n2247_o | n2250_o;
  /* TG68KdotC_Kernel.vhd:1681:103  */
  assign n2252_o = n2251_o & n2240_o;
  /* TG68KdotC_Kernel.vhd:1685:58  */
  assign n2255_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1685:70  */
  assign n2257_o = n2255_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1686:66  */
  assign n2258_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1686:78  */
  assign n2260_o = n2258_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1686:57  */
  assign n2263_o = n2260_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1685:49  */
  assign n2266_o = n2257_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1685:49  */
  assign n2268_o = n2257_o ? n2263_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1691:58  */
  assign n2269_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1691:70  */
  assign n2271_o = n2269_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1691:49  */
  assign n2274_o = n2271_o ? 2'b10 : 2'b00;
  /* TG68KdotC_Kernel.vhd:1696:58  */
  assign n2275_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1696:61  */
  assign n2276_o = ~n2275_o;
  assign n2279_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2280_o = n2305_o ? 1'b1 : n2279_o;
  assign n2281_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2282_o = n2307_o ? 1'b1 : n2281_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2284_o = n2314_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2287_o = n2276_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2289_o = decodeopc & n2276_o;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2291_o = decodeopc & n2276_o;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2292_o = decodeopc & n2276_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2293_o = n2252_o ? n2274_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2295_o = n2252_o ? n2266_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2298_o = n2252_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2301_o = n2252_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2303_o = n2252_o ? n2287_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2305_o = n2289_o & n2252_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2307_o = n2291_o & n2252_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2309_o = n2252_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2311_o = n2252_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2313_o = n2252_o ? n2268_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2314_o = n2292_o & n2252_o;
  /* TG68KdotC_Kernel.vhd:1709:45  */
  assign n2315_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1709:57  */
  assign n2317_o = n2315_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1710:47  */
  assign n2318_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1711:58  */
  assign n2319_o = opcode[11];
  /* TG68KdotC_Kernel.vhd:1712:67  */
  assign n2320_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1712:80  */
  assign n2322_o = n2320_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1713:66  */
  assign n2323_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1713:78  */
  assign n2325_o = n2323_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1712:87  */
  assign n2326_o = n2325_o & n2322_o;
  /* TG68KdotC_Kernel.vhd:1713:96  */
  assign n2327_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1713:108  */
  assign n2329_o = n2327_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1713:125  */
  assign n2330_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1713:137  */
  assign n2332_o = n2330_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1713:116  */
  assign n2333_o = n2329_o | n2332_o;
  /* TG68KdotC_Kernel.vhd:1713:85  */
  assign n2334_o = n2333_o & n2326_o;
  /* TG68KdotC_Kernel.vhd:1714:67  */
  assign n2335_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:1714:86  */
  assign n2336_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1714:98  */
  assign n2338_o = n2336_o == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1714:76  */
  assign n2339_o = n2338_o & n2335_o;
  /* TG68KdotC_Kernel.vhd:1713:145  */
  assign n2340_o = n2334_o | n2339_o;
  /* TG68KdotC_Kernel.vhd:1715:76  */
  assign n2341_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1716:73  */
  assign n2343_o = n2341_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:1717:73  */
  assign n2345_o = n2341_o == 2'b10;
  assign n2346_o = {n2345_o, n2343_o};
  /* TG68KdotC_Kernel.vhd:1715:65  */
  always @*
    case (n2346_o)
      2'b10: n2350_o = 2'b01;
      2'b01: n2350_o = 2'b00;
      default: n2350_o = 2'b10;
    endcase
  /* TG68KdotC_Kernel.vhd:1720:74  */
  assign n2351_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:1720:93  */
  assign n2352_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1720:105  */
  assign n2354_o = n2352_o == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1720:83  */
  assign n2355_o = n2354_o & n2351_o;
  assign n2357_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1721:73  */
  assign n2358_o = decodeopc ? 1'b1 : n2357_o;
  /* TG68KdotC_Kernel.vhd:1721:73  */
  assign n2360_o = decodeopc ? 7'b0111001 : n2180_o;
  assign n2363_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1726:73  */
  assign n2364_o = decodeopc ? 1'b1 : n2363_o;
  assign n2365_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1726:73  */
  assign n2366_o = decodeopc ? 1'b1 : n2365_o;
  /* TG68KdotC_Kernel.vhd:1726:73  */
  assign n2368_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1731:87  */
  assign n2370_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1731:93  */
  assign n2371_o = nextpass & n2370_o;
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2377_o = n2371_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2380_o = n2371_o ? 1'b1 : 1'b0;
  assign n2381_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2382_o = n2371_o ? 1'b1 : n2381_o;
  assign n2383_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2384_o = n2371_o ? 1'b1 : n2383_o;
  assign n2385_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2386_o = n2371_o ? 1'b1 : n2385_o;
  assign n2387_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2388_o = n2371_o ? 1'b1 : n2387_o;
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2390_o = n2371_o ? 7'b0110111 : n2368_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2391_o = n2355_o ? n2026_o : n2377_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2393_o = n2355_o ? 1'b0 : n2380_o;
  assign n2394_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2395_o = n2355_o ? n2394_o : n2382_o;
  assign n2396_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2397_o = n2355_o ? n2396_o : n2364_o;
  assign n2398_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2399_o = n2355_o ? n2398_o : n2384_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2400_o = n2355_o ? n2358_o : n2366_o;
  assign n2401_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2402_o = n2355_o ? n2401_o : n2386_o;
  assign n2403_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2404_o = n2355_o ? n2403_o : n2388_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2405_o = n2355_o ? n2360_o : n2390_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2406_o = n2340_o ? n2350_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2407_o = n2340_o ? n2391_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2409_o = n2340_o ? n2393_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2412_o = n2340_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2415_o = n2340_o ? 1'b0 : 1'b1;
  assign n2416_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2417_o = n2995_o ? n2395_o : n2416_o;
  assign n2418_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2419_o = n2340_o ? n2397_o : n2418_o;
  assign n2420_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2421_o = n2524_o ? n2399_o : n2420_o;
  assign n2422_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2423_o = n2340_o ? n2400_o : n2422_o;
  assign n2424_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2425_o = n3017_o ? n2402_o : n2424_o;
  assign n2426_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2427_o = n3019_o ? n2404_o : n2426_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2428_o = n2340_o ? n2405_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1746:66  */
  assign n2429_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1746:79  */
  assign n2431_o = n2429_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:1747:66  */
  assign n2432_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1747:78  */
  assign n2434_o = n2432_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1746:86  */
  assign n2435_o = n2434_o & n2431_o;
  /* TG68KdotC_Kernel.vhd:1747:95  */
  assign n2436_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1747:107  */
  assign n2438_o = n2436_o != 3'b011;
  /* TG68KdotC_Kernel.vhd:1747:85  */
  assign n2439_o = n2438_o & n2435_o;
  /* TG68KdotC_Kernel.vhd:1747:125  */
  assign n2440_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1747:137  */
  assign n2442_o = n2440_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:1747:115  */
  assign n2443_o = n2442_o & n2439_o;
  /* TG68KdotC_Kernel.vhd:1747:155  */
  assign n2444_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:1747:167  */
  assign n2446_o = n2444_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1747:145  */
  assign n2447_o = n2446_o & n2443_o;
  /* TG68KdotC_Kernel.vhd:1749:83  */
  assign n2449_o = opcode[10:9];
  assign n2452_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1750:65  */
  assign n2453_o = decodeopc ? 1'b1 : n2452_o;
  assign n2454_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2455_o = n2500_o ? 1'b1 : n2454_o;
  /* TG68KdotC_Kernel.vhd:1750:65  */
  assign n2457_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1755:71  */
  assign n2458_o = set[62];
  assign n2461_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2462_o = n2494_o ? 1'b1 : n2461_o;
  assign n2463_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2464_o = n2498_o ? 1'b1 : n2463_o;
  /* TG68KdotC_Kernel.vhd:1759:79  */
  assign n2466_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1759:85  */
  assign n2467_o = nextpass & n2466_o;
  /* TG68KdotC_Kernel.vhd:1762:88  */
  assign n2470_o = exe_datatype != 2'b00;
  /* TG68KdotC_Kernel.vhd:1762:73  */
  assign n2473_o = n2470_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2475_o = n2483_o ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:1759:65  */
  assign n2477_o = n2467_o ? n2473_o : 1'b0;
  assign n2478_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2479_o = n2502_o ? 1'b1 : n2478_o;
  /* TG68KdotC_Kernel.vhd:1759:65  */
  assign n2481_o = n2467_o ? 7'b1000001 : n2457_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2482_o = n2447_o ? n2449_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2483_o = n2467_o & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2486_o = n2447_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2489_o = n2447_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2491_o = n2447_o ? n2477_o : 1'b0;
  assign n2492_o = {1'b1, n2453_o};
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2494_o = n2458_o & n2447_o;
  assign n2495_o = n1909_o[43:42];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2496_o = n2447_o ? n2492_o : n2495_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2498_o = n2458_o & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2500_o = decodeopc & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2502_o = n2467_o & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2503_o = n2447_o ? n2481_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2504_o = n2319_o ? n2406_o : n2482_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2505_o = n2319_o ? n2407_o : n2475_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2507_o = n2319_o ? n2409_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2508_o = n2319_o ? n2412_o : n2486_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2509_o = n2319_o ? n2415_o : n2489_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2511_o = n2319_o ? 1'b0 : n2491_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2513_o = n2340_o & n2319_o;
  assign n2514_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2515_o = n2319_o ? n2514_o : n2462_o;
  assign n2516_o = n2496_o[0];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2517_o = n2319_o ? n2419_o : n2516_o;
  assign n2518_o = n2496_o[1];
  assign n2519_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2520_o = n2319_o ? n2519_o : n2518_o;
  assign n2521_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2522_o = n2319_o ? n2521_o : n2464_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2524_o = n2340_o & n2319_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2525_o = n2319_o ? n2423_o : n2455_o;
  assign n2526_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2527_o = n2319_o ? n2526_o : n2479_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2529_o = n2340_o & n2319_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2531_o = n2340_o & n2319_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2532_o = n2319_o ? n2428_o : n2503_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2533_o = n2979_o ? n2504_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2534_o = n2318_o ? n2505_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2536_o = n2318_o ? n2507_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2538_o = n2318_o ? n2508_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2540_o = n2318_o ? n2509_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2542_o = n2318_o ? n2511_o : 1'b0;
  assign n2543_o = {n2520_o, n2517_o};
  assign n2544_o = {n2421_o, n2522_o};
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2546_o = n2513_o & n2318_o;
  assign n2547_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2548_o = n2997_o ? n2515_o : n2547_o;
  assign n2549_o = n1909_o[43:42];
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2550_o = n2318_o ? n2543_o : n2549_o;
  assign n2551_o = n1909_o[56:55];
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2552_o = n2318_o ? n2544_o : n2551_o;
  assign n2553_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2554_o = n2318_o ? n2525_o : n2553_o;
  assign n2555_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2556_o = n3015_o ? n2527_o : n2555_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2558_o = n2529_o & n2318_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2560_o = n2531_o & n2318_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2561_o = n2318_o ? n2532_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1776:45  */
  assign n2562_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1776:58  */
  assign n2564_o = n2562_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1777:47  */
  assign n2565_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:1777:65  */
  assign n2566_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1777:77  */
  assign n2568_o = n2566_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:1777:55  */
  assign n2569_o = n2568_o & n2565_o;
  /* TG68KdotC_Kernel.vhd:1777:94  */
  assign n2570_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1777:106  */
  assign n2572_o = n2570_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1777:84  */
  assign n2573_o = n2572_o & n2569_o;
  /* TG68KdotC_Kernel.vhd:1777:124  */
  assign n2574_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1777:136  */
  assign n2576_o = n2574_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1777:153  */
  assign n2577_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1777:165  */
  assign n2579_o = n2577_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1777:144  */
  assign n2580_o = n2576_o | n2579_o;
  /* TG68KdotC_Kernel.vhd:1777:113  */
  assign n2581_o = n2580_o & n2573_o;
  /* TG68KdotC_Kernel.vhd:1778:49  */
  assign n2584_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:49  */
  assign n2587_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1777:41  */
  assign n2589_o = n2581_o ? n2584_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1777:41  */
  assign n2591_o = n2581_o ? n2587_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:50  */
  assign n2592_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1791:62  */
  assign n2594_o = n2592_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:1791:79  */
  assign n2595_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1791:91  */
  assign n2597_o = n2595_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1791:69  */
  assign n2598_o = n2597_o & n2594_o;
  /* TG68KdotC_Kernel.vhd:1792:58  */
  assign n2599_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1792:71  */
  assign n2601_o = n2599_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1793:66  */
  assign n2602_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1793:78  */
  assign n2604_o = n2602_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1793:95  */
  assign n2605_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1793:107  */
  assign n2607_o = n2605_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1793:86  */
  assign n2608_o = n2604_o | n2607_o;
  /* TG68KdotC_Kernel.vhd:1793:123  */
  assign n2609_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1793:135  */
  assign n2611_o = n2609_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1793:152  */
  assign n2612_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1793:155  */
  assign n2613_o = ~n2612_o;
  /* TG68KdotC_Kernel.vhd:1793:142  */
  assign n2614_o = n2613_o & n2611_o;
  /* TG68KdotC_Kernel.vhd:1793:113  */
  assign n2615_o = n2608_o | n2614_o;
  /* TG68KdotC_Kernel.vhd:1793:57  */
  assign n2619_o = n2615_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1793:57  */
  assign n2622_o = n2615_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1793:57  */
  assign n2624_o = n2615_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1792:49  */
  assign n2626_o = n2601_o ? n2619_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1792:49  */
  assign n2628_o = n2601_o ? n2622_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1792:49  */
  assign n2630_o = n2601_o ? n2624_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1800:58  */
  assign n2631_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1800:71  */
  assign n2633_o = n2631_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1801:66  */
  assign n2634_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1801:78  */
  assign n2636_o = n2634_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1801:95  */
  assign n2637_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1801:107  */
  assign n2639_o = n2637_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1801:86  */
  assign n2640_o = n2636_o | n2639_o;
  /* TG68KdotC_Kernel.vhd:1801:123  */
  assign n2641_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1801:135  */
  assign n2643_o = n2641_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1801:152  */
  assign n2644_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1801:155  */
  assign n2645_o = ~n2644_o;
  /* TG68KdotC_Kernel.vhd:1801:142  */
  assign n2646_o = n2645_o & n2643_o;
  /* TG68KdotC_Kernel.vhd:1801:113  */
  assign n2647_o = n2640_o | n2646_o;
  /* TG68KdotC_Kernel.vhd:1801:57  */
  assign n2650_o = n2647_o ? n2626_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1801:57  */
  assign n2652_o = n2647_o ? n2628_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1801:57  */
  assign n2654_o = n2647_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1800:49  */
  assign n2655_o = n2633_o ? n2650_o : n2626_o;
  /* TG68KdotC_Kernel.vhd:1800:49  */
  assign n2656_o = n2633_o ? n2652_o : n2628_o;
  /* TG68KdotC_Kernel.vhd:1800:49  */
  assign n2658_o = n2633_o ? n2654_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1808:58  */
  assign n2659_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1808:71  */
  assign n2661_o = n2659_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1808:87  */
  assign n2662_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1808:100  */
  assign n2664_o = n2662_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1808:78  */
  assign n2665_o = n2661_o | n2664_o;
  /* TG68KdotC_Kernel.vhd:1809:66  */
  assign n2666_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1809:78  */
  assign n2668_o = n2666_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1809:95  */
  assign n2669_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1809:107  */
  assign n2671_o = n2669_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1809:86  */
  assign n2672_o = n2668_o | n2671_o;
  /* TG68KdotC_Kernel.vhd:1809:57  */
  assign n2675_o = n2672_o ? n2655_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1809:57  */
  assign n2677_o = n2672_o ? n2656_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1809:57  */
  assign n2679_o = n2672_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1808:49  */
  assign n2680_o = n2665_o ? n2675_o : n2655_o;
  /* TG68KdotC_Kernel.vhd:1808:49  */
  assign n2681_o = n2665_o ? n2677_o : n2656_o;
  /* TG68KdotC_Kernel.vhd:1808:49  */
  assign n2683_o = n2665_o ? n2679_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1816:58  */
  assign n2684_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1816:71  */
  assign n2686_o = n2684_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:1817:66  */
  assign n2687_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1817:78  */
  assign n2689_o = n2687_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1817:95  */
  assign n2690_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1817:107  */
  assign n2692_o = n2690_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1817:86  */
  assign n2693_o = n2689_o | n2692_o;
  /* TG68KdotC_Kernel.vhd:1817:123  */
  assign n2694_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1817:135  */
  assign n2696_o = n2694_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1817:152  */
  assign n2697_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1817:155  */
  assign n2698_o = ~n2697_o;
  /* TG68KdotC_Kernel.vhd:1817:142  */
  assign n2699_o = n2698_o & n2696_o;
  /* TG68KdotC_Kernel.vhd:1817:113  */
  assign n2700_o = n2693_o | n2699_o;
  /* TG68KdotC_Kernel.vhd:1817:57  */
  assign n2703_o = n2700_o ? n2680_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1817:57  */
  assign n2705_o = n2700_o ? n2681_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1817:57  */
  assign n2707_o = n2700_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1816:49  */
  assign n2708_o = n2686_o ? n2703_o : n2680_o;
  /* TG68KdotC_Kernel.vhd:1816:49  */
  assign n2709_o = n2686_o ? n2705_o : n2681_o;
  /* TG68KdotC_Kernel.vhd:1816:49  */
  assign n2711_o = n2686_o ? n2707_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1824:58  */
  assign n2712_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1824:71  */
  assign n2714_o = n2712_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:1825:66  */
  assign n2715_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1825:78  */
  assign n2717_o = n2715_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1825:95  */
  assign n2718_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:1825:98  */
  assign n2719_o = ~n2718_o;
  /* TG68KdotC_Kernel.vhd:1825:86  */
  assign n2720_o = n2717_o | n2719_o;
  /* TG68KdotC_Kernel.vhd:1825:57  */
  assign n2723_o = n2720_o ? n2708_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1825:57  */
  assign n2725_o = n2720_o ? n2709_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1825:57  */
  assign n2727_o = n2720_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1824:49  */
  assign n2728_o = n2714_o ? n2723_o : n2708_o;
  /* TG68KdotC_Kernel.vhd:1824:49  */
  assign n2729_o = n2714_o ? n2725_o : n2709_o;
  /* TG68KdotC_Kernel.vhd:1824:49  */
  assign n2731_o = n2714_o ? n2727_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1832:61  */
  assign n2732_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1832:80  */
  assign n2733_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1832:69  */
  assign n2734_o = n2732_o | n2733_o;
  /* TG68KdotC_Kernel.vhd:1832:100  */
  assign n2735_o = set_exec[3];
  /* TG68KdotC_Kernel.vhd:1832:89  */
  assign n2736_o = n2734_o | n2735_o;
  /* TG68KdotC_Kernel.vhd:1832:120  */
  assign n2737_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1832:109  */
  assign n2738_o = n2736_o | n2737_o;
  /* TG68KdotC_Kernel.vhd:1832:140  */
  assign n2739_o = set_exec[8];
  /* TG68KdotC_Kernel.vhd:1832:129  */
  assign n2740_o = n2738_o | n2739_o;
  /* TG68KdotC_Kernel.vhd:1833:66  */
  assign n2741_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1833:69  */
  assign n2742_o = ~n2741_o;
  /* TG68KdotC_Kernel.vhd:1833:84  */
  assign n2743_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1833:96  */
  assign n2745_o = n2743_o == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1833:74  */
  assign n2746_o = n2745_o & n2742_o;
  /* TG68KdotC_Kernel.vhd:1833:119  */
  assign n2747_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1833:139  */
  assign n2748_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1833:128  */
  assign n2749_o = n2747_o | n2748_o;
  /* TG68KdotC_Kernel.vhd:1833:158  */
  assign n2750_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1833:147  */
  assign n2751_o = n2749_o | n2750_o;
  /* TG68KdotC_Kernel.vhd:1833:106  */
  assign n2752_o = n2751_o & n2746_o;
  /* TG68KdotC_Kernel.vhd:1834:92  */
  assign n2753_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:1834:82  */
  assign n2754_o = n2753_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1834:107  */
  assign n2755_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1834:97  */
  assign n2756_o = n2755_o & n2754_o;
  /* TG68KdotC_Kernel.vhd:1840:90  */
  assign n2758_o = opcode[6];
  assign n2760_o = n1909_o[52];
  /* TG68KdotC_Kernel.vhd:1840:81  */
  assign n2761_o = n2758_o ? 1'b1 : n2760_o;
  /* TG68KdotC_Kernel.vhd:1844:104  */
  assign n2763_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1845:104  */
  assign n2764_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1846:103  */
  assign n2765_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2767_o = decodeopc ? 2'b01 : n2026_o;
  assign n2768_o = {n2765_o, n2764_o, n2763_o};
  assign n2769_o = {n2761_o, 1'b1};
  assign n2770_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2771_o = decodeopc ? n2768_o : n2770_o;
  assign n2772_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2773_o = decodeopc ? n2769_o : n2772_o;
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2775_o = decodeopc ? 7'b0011000 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2776_o = n2756_o ? n2026_o : n2767_o;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2779_o = n2756_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2781_o = n2756_o ? 1'b1 : n2729_o;
  assign n2782_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2783_o = n2756_o ? n2782_o : n2771_o;
  assign n2784_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2785_o = n2756_o ? n2784_o : 1'b1;
  assign n2786_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2787_o = n2756_o ? n2786_o : n2773_o;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2788_o = n2756_o ? n2180_o : n2775_o;
  /* TG68KdotC_Kernel.vhd:1851:69  */
  assign n2789_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1851:72  */
  assign n2790_o = ~n2789_o;
  /* TG68KdotC_Kernel.vhd:1851:86  */
  assign n2791_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1851:98  */
  assign n2793_o = n2791_o != 6'b111100;
  /* TG68KdotC_Kernel.vhd:1851:77  */
  assign n2794_o = n2790_o | n2793_o;
  /* TG68KdotC_Kernel.vhd:1851:121  */
  assign n2795_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1851:141  */
  assign n2796_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1851:130  */
  assign n2797_o = n2795_o | n2796_o;
  /* TG68KdotC_Kernel.vhd:1851:160  */
  assign n2798_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1851:149  */
  assign n2799_o = n2797_o | n2798_o;
  /* TG68KdotC_Kernel.vhd:1851:169  */
  assign n2800_o = ~n2799_o;
  /* TG68KdotC_Kernel.vhd:1851:109  */
  assign n2801_o = n2794_o | n2800_o;
  /* TG68KdotC_Kernel.vhd:1857:84  */
  assign n2805_o = datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2807_o = n2856_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2809_o = n2845_o ? 1'b1 : n2154_o;
  assign n2810_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2811_o = n2851_o ? 1'b1 : n2810_o;
  assign n2812_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2813_o = n2855_o ? 1'b1 : n2812_o;
  /* TG68KdotC_Kernel.vhd:1852:65  */
  assign n2814_o = n2805_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2816_o = n2861_o ? 7'b0011101 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1861:74  */
  assign n2817_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1861:86  */
  assign n2819_o = n2817_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1861:65  */
  assign n2822_o = n2819_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1864:74  */
  assign n2823_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1864:87  */
  assign n2825_o = n2823_o != 3'b110;
  /* TG68KdotC_Kernel.vhd:1865:82  */
  assign n2826_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1865:94  */
  assign n2828_o = n2826_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1865:73  */
  assign n2831_o = n2828_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1864:65  */
  assign n2834_o = n2825_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1864:65  */
  assign n2836_o = n2825_o ? n2831_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1870:74  */
  assign n2837_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1870:87  */
  assign n2839_o = n2837_o == 2'b10;
  assign n2841_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2842_o = n2853_o ? 1'b1 : n2841_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2844_o = n2801_o ? n2834_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2845_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2847_o = n2801_o ? n2728_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2849_o = n2801_o ? n2729_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2851_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2853_o = n2839_o & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2855_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2856_o = n2814_o & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2858_o = n2801_o ? n2822_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2860_o = n2801_o ? n2836_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2861_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2862_o = n2916_o ? n2776_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2864_o = n2752_o ? 1'b0 : n2844_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2865_o = n2752_o ? n2154_o : n2809_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2866_o = n2752_o ? n2728_o : n2847_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2868_o = n2752_o ? n2779_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2869_o = n2752_o ? n2781_o : n2849_o;
  assign n2870_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2871_o = n2927_o ? n2783_o : n2870_o;
  assign n2872_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2873_o = n2752_o ? n2872_o : n2811_o;
  assign n2874_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2875_o = n2931_o ? n2785_o : n2874_o;
  assign n2876_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2877_o = n2933_o ? n2787_o : n2876_o;
  assign n2878_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2879_o = n2752_o ? n2878_o : n2842_o;
  assign n2880_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2881_o = n2752_o ? n2880_o : n2813_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2882_o = n2752_o ? n2171_o : n2807_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2884_o = n2752_o ? 1'b0 : n2858_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2886_o = n2752_o ? 1'b0 : n2860_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2887_o = n2752_o ? n2788_o : n2816_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2888_o = n2752_o & n2740_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2890_o = n2740_o ? n2864_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2891_o = n2919_o ? n2865_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2893_o = n2740_o ? n2866_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2895_o = n2740_o ? n2868_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2897_o = n2740_o ? n2869_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2899_o = n2752_o & n2740_o;
  assign n2900_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2901_o = n2929_o ? n2873_o : n2900_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2903_o = n2752_o & n2740_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2905_o = n2752_o & n2740_o;
  assign n2906_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2907_o = n2935_o ? n2879_o : n2906_o;
  assign n2908_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2909_o = n2937_o ? n2881_o : n2908_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2910_o = n2938_o ? n2882_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2912_o = n2740_o ? n2884_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2914_o = n2740_o ? n2886_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2915_o = n2948_o ? n2887_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2916_o = n2888_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2918_o = n2598_o ? n2890_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2919_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2921_o = n2598_o ? n2893_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2923_o = n2598_o ? n2895_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2925_o = n2598_o ? n2897_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2927_o = n2899_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2929_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2931_o = n2903_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2933_o = n2905_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2935_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2937_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2938_o = n2740_o & n2598_o;
  assign n2939_o = {n2731_o, n2711_o, n2658_o, n2630_o};
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2941_o = n2598_o ? n2683_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2943_o = n2598_o ? n2939_o : 4'b0000;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2945_o = n2598_o ? n2912_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2947_o = n2598_o ? n2914_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2948_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2949_o = n2564_o ? n2026_o : n2862_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2951_o = n2564_o ? 1'b0 : n2918_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2952_o = n2564_o ? n2154_o : n2891_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2953_o = n2564_o ? n2589_o : n2921_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2954_o = n2564_o ? n2591_o : n2923_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2956_o = n2564_o ? 1'b1 : n2925_o;
  assign n2957_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2958_o = n2564_o ? n2957_o : n2871_o;
  assign n2959_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2960_o = n2564_o ? n2959_o : n2901_o;
  assign n2961_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2962_o = n2564_o ? n2961_o : n2875_o;
  assign n2963_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2964_o = n2564_o ? n2963_o : n2877_o;
  assign n2965_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2966_o = n2564_o ? n2965_o : n2907_o;
  assign n2967_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2968_o = n2564_o ? n2967_o : n2909_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2969_o = n2564_o ? n2171_o : n2910_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2971_o = n2564_o ? 1'b0 : n2941_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2973_o = n2564_o ? 4'b0000 : n2943_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2975_o = n2564_o ? 1'b0 : n2945_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2977_o = n2564_o ? 1'b0 : n2947_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2978_o = n2564_o ? n2180_o : n2915_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2979_o = n2318_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2980_o = n2317_o ? n2534_o : n2949_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2982_o = n2317_o ? 1'b0 : n2951_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2984_o = n2317_o ? n2536_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2985_o = n2317_o ? n2154_o : n2952_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2986_o = n2317_o ? n2538_o : n2953_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2988_o = n2317_o ? 1'b0 : n2954_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2989_o = n2317_o ? n2540_o : n2956_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2991_o = n2317_o ? n2542_o : 1'b0;
  assign n2992_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2993_o = n2317_o ? n2992_o : n2958_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2995_o = n2546_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2997_o = n2318_o & n2317_o;
  assign n2998_o = n2550_o[0];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2999_o = n2317_o ? n2998_o : n2960_o;
  assign n3000_o = n2550_o[1];
  assign n3001_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3002_o = n2317_o ? n3000_o : n3001_o;
  assign n3003_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3004_o = n2317_o ? n3003_o : n2962_o;
  assign n3005_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3006_o = n2317_o ? n3005_o : n2964_o;
  assign n3007_o = n2552_o[0];
  assign n3008_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3009_o = n2317_o ? n3007_o : n3008_o;
  assign n3010_o = n2552_o[1];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3011_o = n2317_o ? n3010_o : n2966_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3012_o = n2317_o ? n2554_o : n2968_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3013_o = n2317_o ? n2171_o : n2969_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3015_o = n2318_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3017_o = n2558_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3019_o = n2560_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3021_o = n2317_o ? 1'b0 : n2971_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3023_o = n2317_o ? 4'b0000 : n2973_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3025_o = n2317_o ? 1'b0 : n2975_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3027_o = n2317_o ? 1'b0 : n2977_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3028_o = n2317_o ? n2561_o : n2978_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3029_o = n2222_o ? n2293_o : n2533_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3030_o = n2222_o ? n2026_o : n2980_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3031_o = n2222_o ? n2295_o : n2982_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3033_o = n2222_o ? 1'b0 : n2984_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3034_o = n2222_o ? n2154_o : n2985_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3035_o = n2222_o ? n2298_o : n2986_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3037_o = n2222_o ? 1'b0 : n2988_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3038_o = n2222_o ? n2301_o : n2989_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3040_o = n2222_o ? n2303_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3042_o = n2222_o ? 1'b0 : n2991_o;
  assign n3043_o = {n3002_o, n2999_o};
  assign n3044_o = {n3011_o, n3009_o};
  assign n3045_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3046_o = n2222_o ? n3045_o : n2993_o;
  assign n3047_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3048_o = n2222_o ? n3047_o : n2417_o;
  assign n3049_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3050_o = n2222_o ? n3049_o : n2548_o;
  assign n3051_o = n3043_o[0];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3052_o = n2222_o ? n2280_o : n3051_o;
  assign n3053_o = n3043_o[1];
  assign n3054_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3055_o = n2222_o ? n3054_o : n3053_o;
  assign n3056_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3057_o = n2222_o ? n3056_o : n3004_o;
  assign n3058_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3059_o = n2222_o ? n3058_o : n3006_o;
  assign n3060_o = n1909_o[56:55];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3061_o = n2222_o ? n3060_o : n3044_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3062_o = n2222_o ? n2282_o : n3012_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3063_o = n2222_o ? n2171_o : n3013_o;
  assign n3064_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3065_o = n2222_o ? n3064_o : n2556_o;
  assign n3066_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3067_o = n2222_o ? n3066_o : n2425_o;
  assign n3068_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3069_o = n2222_o ? n3068_o : n2427_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3071_o = n2222_o ? 1'b0 : n3021_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3073_o = n2222_o ? 4'b0000 : n3023_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3075_o = n2222_o ? n2309_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3076_o = n2222_o ? n2311_o : n3025_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3077_o = n2222_o ? n2313_o : n3027_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3078_o = n2222_o ? n2284_o : n3028_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3080_o = n2190_o ? 2'b00 : n3029_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3081_o = n2190_o ? n2026_o : n3030_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3083_o = n2190_o ? 1'b0 : n3031_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3085_o = n2190_o ? 1'b0 : n3033_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3087_o = n2190_o ? n2217_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3088_o = n2190_o ? n2210_o : n3034_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3090_o = n2190_o ? 1'b0 : n3035_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3092_o = n2190_o ? 1'b0 : n3037_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3094_o = n2190_o ? 1'b0 : n3038_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3096_o = n2190_o ? 1'b0 : n3040_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3098_o = n2190_o ? 1'b0 : n3042_o;
  assign n3099_o = {n3055_o, n3052_o};
  assign n3100_o = {1'b1, 1'b1};
  assign n3101_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3102_o = n2190_o ? n3101_o : n3046_o;
  assign n3103_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3104_o = n2190_o ? n3103_o : n3048_o;
  assign n3105_o = n1909_o[37];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3106_o = n2190_o ? n2206_o : n3105_o;
  assign n3107_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3108_o = n2190_o ? n3107_o : n3050_o;
  assign n3109_o = n1909_o[43:42];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3110_o = n2190_o ? n3109_o : n3099_o;
  assign n3111_o = n3100_o[0];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3112_o = n2190_o ? n3111_o : n3057_o;
  assign n3113_o = n3100_o[1];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3114_o = n2190_o ? n3113_o : n2168_o;
  assign n3115_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3116_o = n2190_o ? n3115_o : n3059_o;
  assign n3117_o = n1909_o[56:55];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3118_o = n2190_o ? n3117_o : n3061_o;
  assign n3119_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3120_o = n2190_o ? n3119_o : n3062_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3121_o = n2190_o ? n2171_o : n3063_o;
  assign n3122_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3123_o = n2190_o ? n3122_o : n3065_o;
  assign n3124_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3125_o = n2190_o ? n3124_o : n3067_o;
  assign n3126_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3127_o = n2190_o ? n3126_o : n3069_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3129_o = n2190_o ? n2201_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3131_o = n2190_o ? 1'b0 : n3071_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3133_o = n2190_o ? 4'b0000 : n3073_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3135_o = n2190_o ? 1'b0 : n3075_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3137_o = n2190_o ? 1'b0 : n3076_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3138_o = n2190_o ? n2203_o : n3077_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3139_o = n2190_o ? n2214_o : n3078_o;
  /* TG68KdotC_Kernel.vhd:1655:25  */
  assign n3141_o = n2185_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:1890:44  */
  assign n3142_o = opcode[11:10];
  /* TG68KdotC_Kernel.vhd:1890:58  */
  assign n3144_o = n3142_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1890:73  */
  assign n3145_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1890:85  */
  assign n3147_o = n3145_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1890:64  */
  assign n3148_o = n3144_o | n3147_o;
  /* TG68KdotC_Kernel.vhd:1891:43  */
  assign n3149_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:1891:55  */
  assign n3151_o = n3149_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1891:73  */
  assign n3152_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:1891:85  */
  assign n3154_o = n3152_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1891:64  */
  assign n3155_o = n3151_o | n3154_o;
  /* TG68KdotC_Kernel.vhd:1890:94  */
  assign n3156_o = n3155_o & n3148_o;
  /* TG68KdotC_Kernel.vhd:1892:43  */
  assign n3157_o = opcode[13];
  /* TG68KdotC_Kernel.vhd:1892:62  */
  assign n3158_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1892:74  */
  assign n3160_o = n3158_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1892:92  */
  assign n3161_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1892:104  */
  assign n3163_o = n3161_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1892:82  */
  assign n3164_o = n3163_o & n3160_o;
  /* TG68KdotC_Kernel.vhd:1892:52  */
  assign n3165_o = n3157_o | n3164_o;
  /* TG68KdotC_Kernel.vhd:1891:92  */
  assign n3166_o = n3165_o & n3156_o;
  /* TG68KdotC_Kernel.vhd:1895:50  */
  assign n3168_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1895:62  */
  assign n3170_o = n3168_o == 3'b001;
  assign n3172_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1895:41  */
  assign n3173_o = n3170_o ? 1'b1 : n3172_o;
  /* TG68KdotC_Kernel.vhd:1898:50  */
  assign n3174_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1898:62  */
  assign n3176_o = n3174_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1899:58  */
  assign n3177_o = opcode[8:7];
  /* TG68KdotC_Kernel.vhd:1899:70  */
  assign n3179_o = n3177_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1899:49  */
  assign n3182_o = n3179_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1898:41  */
  assign n3184_o = n3176_o ? n3182_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1903:52  */
  assign n3185_o = opcode[13:12];
  /* TG68KdotC_Kernel.vhd:1904:49  */
  assign n3187_o = n3185_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:1905:49  */
  assign n3189_o = n3185_o == 2'b10;
  assign n3190_o = {n3189_o, n3187_o};
  /* TG68KdotC_Kernel.vhd:1903:41  */
  always @*
    case (n3190_o)
      2'b10: n3194_o = 2'b10;
      2'b01: n3194_o = 2'b00;
      default: n3194_o = 2'b01;
    endcase
  /* TG68KdotC_Kernel.vhd:1909:50  */
  assign n3195_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:1909:41  */
  assign n3198_o = n3195_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1913:66  */
  assign n3199_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1913:78  */
  assign n3201_o = n3199_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1913:57  */
  assign n3202_o = nextpass | n3201_o;
  /* TG68KdotC_Kernel.vhd:1915:58  */
  assign n3203_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1915:70  */
  assign n3205_o = n3203_o != 3'b000;
  /* TG68KdotC_Kernel.vhd:1915:49  */
  assign n3208_o = n3205_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1913:41  */
  assign n3210_o = n3202_o ? n3208_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1913:41  */
  assign n3213_o = n3202_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1920:55  */
  assign n3215_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1920:89  */
  assign n3216_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1920:101  */
  assign n3218_o = n3216_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1920:107  */
  assign n3219_o = decodeopc & n3218_o;
  /* TG68KdotC_Kernel.vhd:1920:79  */
  assign n3220_o = nextpass | n3219_o;
  /* TG68KdotC_Kernel.vhd:1920:61  */
  assign n3221_o = n3220_o & n3215_o;
  /* TG68KdotC_Kernel.vhd:1921:60  */
  assign n3222_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1922:57  */
  assign n3225_o = n3222_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1922:67  */
  assign n3227_o = n3222_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1922:67  */
  assign n3228_o = n3225_o | n3227_o;
  /* TG68KdotC_Kernel.vhd:1925:74  */
  assign n3229_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1927:82  */
  assign n3231_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1927:95  */
  assign n3233_o = n3231_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1925:65  */
  assign n3235_o = n3240_o ? 1'b1 : n2168_o;
  assign n3236_o = n2162_o[0];
  assign n3237_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3238_o = n2037_o ? n3236_o : n3237_o;
  /* TG68KdotC_Kernel.vhd:1925:65  */
  assign n3239_o = n3229_o ? 1'b1 : n3238_o;
  /* TG68KdotC_Kernel.vhd:1925:65  */
  assign n3240_o = n3233_o & n3229_o;
  /* TG68KdotC_Kernel.vhd:1931:74  */
  assign n3241_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1933:82  */
  assign n3243_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1933:95  */
  assign n3245_o = n3243_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1931:65  */
  assign n3247_o = n3252_o ? 1'b1 : n3235_o;
  assign n3248_o = n2162_o[1];
  assign n3249_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3250_o = n2037_o ? n3248_o : n3249_o;
  /* TG68KdotC_Kernel.vhd:1931:65  */
  assign n3251_o = n3241_o ? 1'b1 : n3250_o;
  /* TG68KdotC_Kernel.vhd:1931:65  */
  assign n3252_o = n3245_o & n3241_o;
  /* TG68KdotC_Kernel.vhd:1939:76  */
  assign n3253_o = ~nextpass;
  assign n3255_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1939:65  */
  assign n3256_o = n3253_o ? 1'b1 : n3255_o;
  /* TG68KdotC_Kernel.vhd:1924:57  */
  assign n3258_o = n3222_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1924:67  */
  assign n3260_o = n3222_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1924:67  */
  assign n3261_o = n3258_o | n3260_o;
  /* TG68KdotC_Kernel.vhd:1924:73  */
  assign n3263_o = n3222_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1924:73  */
  assign n3264_o = n3261_o | n3263_o;
  /* TG68KdotC_Kernel.vhd:1942:57  */
  assign n3266_o = n3222_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:1945:57  */
  assign n3268_o = n3222_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:1949:76  */
  assign n3269_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1950:73  */
  assign n3271_o = n3269_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1952:73  */
  assign n3274_o = n3269_o == 3'b001;
  assign n3275_o = {n3274_o, n3271_o};
  /* TG68KdotC_Kernel.vhd:1949:65  */
  always @*
    case (n3275_o)
      2'b10: n3276_o = 1'b1;
      2'b01: n3276_o = n2171_o;
      default: n3276_o = n2171_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1949:65  */
  always @*
    case (n3275_o)
      2'b10: n3279_o = 7'b0000011;
      2'b01: n3279_o = 7'b0000011;
      default: n3279_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1948:57  */
  assign n3281_o = n3222_o == 3'b111;
  assign n3282_o = {n3281_o, n3268_o, n3266_o, n3264_o, n3228_o};
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3284_o = n2026_o;
      5'b01000: n3284_o = n2026_o;
      5'b00100: n3284_o = n2026_o;
      5'b00010: n3284_o = 2'b11;
      5'b00001: n3284_o = n2026_o;
      default: n3284_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3286_o = n2151_o;
      5'b01000: n3286_o = 1'b1;
      5'b00100: n3286_o = n2151_o;
      5'b00010: n3286_o = n2151_o;
      5'b00001: n3286_o = n2151_o;
      default: n3286_o = n2151_o;
    endcase
  assign n3287_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3288_o = n3287_o;
      5'b01000: n3288_o = n3287_o;
      5'b00100: n3288_o = n3287_o;
      5'b00010: n3288_o = n3256_o;
      5'b00001: n3288_o = n3287_o;
      default: n3288_o = n3287_o;
    endcase
  assign n3289_o = n2162_o[0];
  assign n3290_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3291_o = n2037_o ? n3289_o : n3290_o;
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3292_o = n3291_o;
      5'b01000: n3292_o = n3291_o;
      5'b00100: n3292_o = n3291_o;
      5'b00010: n3292_o = n3239_o;
      5'b00001: n3292_o = n3291_o;
      default: n3292_o = n3291_o;
    endcase
  assign n3293_o = n2162_o[1];
  assign n3294_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3295_o = n2037_o ? n3293_o : n3294_o;
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3296_o = n3295_o;
      5'b01000: n3296_o = n3295_o;
      5'b00100: n3296_o = n3295_o;
      5'b00010: n3296_o = n3251_o;
      5'b00001: n3296_o = n3295_o;
      default: n3296_o = n3295_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3297_o = n2168_o;
      5'b01000: n3297_o = n2168_o;
      5'b00100: n3297_o = n2168_o;
      5'b00010: n3297_o = n3247_o;
      5'b00001: n3297_o = n2168_o;
      default: n3297_o = n2168_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3298_o = n3276_o;
      5'b01000: n3298_o = n2171_o;
      5'b00100: n3298_o = n2171_o;
      5'b00010: n3298_o = n2171_o;
      5'b00001: n3298_o = n2171_o;
      default: n3298_o = n2171_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3299_o = n3184_o;
      5'b01000: n3299_o = n3184_o;
      5'b00100: n3299_o = n3184_o;
      5'b00010: n3299_o = n3184_o;
      5'b00001: n3299_o = 1'b1;
      default: n3299_o = n3184_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3303_o = n3279_o;
      5'b01000: n3303_o = 7'b0010011;
      5'b00100: n3303_o = 7'b0000111;
      5'b00010: n3303_o = 7'b0000001;
      5'b00001: n3303_o = n2180_o;
      default: n3303_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3304_o = n3315_o ? n3284_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3305_o = n3316_o ? n3286_o : n2151_o;
  assign n3306_o = {n3296_o, n3292_o};
  assign n3307_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3308_o = n3337_o ? n3288_o : n3307_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3309_o = n3338_o ? n3306_o : n2166_o;
  /* TG68KdotC_Kernel.vhd:1920:41  */
  assign n3310_o = n3221_o ? n3297_o : n2168_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3311_o = n3342_o ? n3298_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:1920:41  */
  assign n3312_o = n3221_o ? n3299_o : n3184_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3313_o = n3347_o ? n3303_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3314_o = n3166_o ? n3194_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3315_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3316_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3318_o = n3166_o ? n3198_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3321_o = n3166_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3323_o = n3166_o ? n3210_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3325_o = n3166_o ? n3213_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3328_o = n3166_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3331_o = n3166_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3334_o = n3166_o ? 1'b1 : 1'b0;
  assign n3335_o = {n3310_o, n3173_o};
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3337_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3338_o = n3221_o & n3166_o;
  assign n3339_o = n1909_o[49];
  assign n3340_o = {n2168_o, n3339_o};
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3341_o = n3166_o ? n3335_o : n3340_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3342_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3344_o = n3166_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3346_o = n3166_o ? n3312_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3347_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1889:25  */
  assign n3349_o = n2185_o == 4'b0001;
  /* TG68KdotC_Kernel.vhd:1889:36  */
  assign n3351_o = n2185_o == 4'b0010;
  /* TG68KdotC_Kernel.vhd:1889:36  */
  assign n3352_o = n3349_o | n3351_o;
  /* TG68KdotC_Kernel.vhd:1889:43  */
  assign n3354_o = n2185_o == 4'b0011;
  /* TG68KdotC_Kernel.vhd:1889:43  */
  assign n3355_o = n3352_o | n3354_o;
  /* TG68KdotC_Kernel.vhd:1966:42  */
  assign n3356_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1967:50  */
  assign n3357_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1968:58  */
  assign n3358_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1968:71  */
  assign n3360_o = n3358_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1968:88  */
  assign n3361_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1968:100  */
  assign n3363_o = n3361_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1968:78  */
  assign n3364_o = n3363_o & n3360_o;
  /* TG68KdotC_Kernel.vhd:1969:66  */
  assign n3365_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1969:81  */
  assign n3366_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1969:74  */
  assign n3367_o = n3366_o & n3365_o;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3374_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3377_o = n3367_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3380_o = n3367_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3382_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3384_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3386_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3388_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:66  */
  assign n3389_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1981:67  */
  assign n3390_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:1981:84  */
  assign n3391_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:1981:96  */
  assign n3393_o = n3391_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:1981:75  */
  assign n3394_o = n3390_o | n3393_o;
  /* TG68KdotC_Kernel.vhd:1980:74  */
  assign n3395_o = n3394_o & n3389_o;
  /* TG68KdotC_Kernel.vhd:1982:66  */
  assign n3396_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1982:78  */
  assign n3398_o = n3396_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:1981:103  */
  assign n3399_o = n3398_o & n3395_o;
  /* TG68KdotC_Kernel.vhd:1982:96  */
  assign n3400_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:1982:108  */
  assign n3402_o = n3400_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1982:86  */
  assign n3403_o = n3402_o & n3399_o;
  /* TG68KdotC_Kernel.vhd:1989:74  */
  assign n3407_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1989:86  */
  assign n3409_o = n3407_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1989:65  */
  assign n3412_o = n3409_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1989:65  */
  assign n3415_o = n3409_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1989:65  */
  assign n3418_o = n3409_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1995:71  */
  assign n3419_o = set[62];
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3421_o = n3428_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3423_o = n3442_o ? 1'b1 : n2154_o;
  /* TG68KdotC_Kernel.vhd:1999:65  */
  assign n3425_o = setexecopc ? 1'b1 : n3412_o;
  /* TG68KdotC_Kernel.vhd:1999:65  */
  assign n3427_o = setexecopc ? 1'b1 : n3415_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3428_o = n3419_o & n3403_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3431_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3434_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3437_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3439_o = n3403_o ? n3425_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3441_o = n3403_o ? n3427_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3442_o = n3419_o & n3403_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3445_o = n3403_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3448_o = n3403_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3450_o = n3403_o ? n3418_o : 1'b0;
  assign n3451_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3452_o = n3403_o ? 1'b1 : n3451_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3454_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3456_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3457_o = n3364_o ? n2026_o : n3421_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3459_o = n3364_o ? 1'b0 : n3431_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3461_o = n3364_o ? 1'b0 : n3434_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3462_o = n3364_o ? n3374_o : n3437_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3464_o = n3364_o ? 1'b0 : n3439_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3466_o = n3364_o ? 1'b0 : n3441_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3467_o = n3364_o ? n2154_o : n3423_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3468_o = n3364_o ? n3377_o : n3445_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3469_o = n3364_o ? n3380_o : n3448_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3471_o = n3364_o ? 1'b0 : n3450_o;
  assign n3472_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3473_o = n3364_o ? n3472_o : n3452_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3474_o = n3364_o ? n3382_o : n3454_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3476_o = n3364_o ? n3384_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3477_o = n3364_o ? n3386_o : n3456_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3479_o = n3364_o ? n3388_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:58  */
  assign n3480_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2009:70  */
  assign n3482_o = n3480_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2010:59  */
  assign n3483_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2010:71  */
  assign n3485_o = n3483_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2010:89  */
  assign n3486_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2010:101  */
  assign n3488_o = n3486_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2010:80  */
  assign n3489_o = n3485_o | n3488_o;
  /* TG68KdotC_Kernel.vhd:2009:78  */
  assign n3490_o = n3489_o & n3482_o;
  /* TG68KdotC_Kernel.vhd:2011:66  */
  assign n3491_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2014:74  */
  assign n3493_o = c_out[1];
  /* TG68KdotC_Kernel.vhd:2014:77  */
  assign n3494_o = ~n3493_o;
  /* TG68KdotC_Kernel.vhd:2014:91  */
  assign n3495_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:2014:82  */
  assign n3496_o = n3494_o | n3495_o;
  /* TG68KdotC_Kernel.vhd:2014:109  */
  assign n3497_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:2014:100  */
  assign n3498_o = n3496_o | n3497_o;
  /* TG68KdotC_Kernel.vhd:2014:127  */
  assign n3499_o = exec[31];
  /* TG68KdotC_Kernel.vhd:2014:119  */
  assign n3500_o = n3499_o & n3498_o;
  /* TG68KdotC_Kernel.vhd:2014:65  */
  assign n3503_o = n3500_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2017:66  */
  assign n3504_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2020:74  */
  assign n3506_o = c_out[2];
  /* TG68KdotC_Kernel.vhd:2020:77  */
  assign n3507_o = ~n3506_o;
  /* TG68KdotC_Kernel.vhd:2020:91  */
  assign n3508_o = op1out[31];
  /* TG68KdotC_Kernel.vhd:2020:82  */
  assign n3509_o = n3507_o | n3508_o;
  /* TG68KdotC_Kernel.vhd:2020:109  */
  assign n3510_o = op2out[31];
  /* TG68KdotC_Kernel.vhd:2020:100  */
  assign n3511_o = n3509_o | n3510_o;
  /* TG68KdotC_Kernel.vhd:2020:127  */
  assign n3512_o = exec[31];
  /* TG68KdotC_Kernel.vhd:2020:119  */
  assign n3513_o = n3512_o & n3511_o;
  /* TG68KdotC_Kernel.vhd:2020:65  */
  assign n3516_o = n3513_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3518_o = n3504_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3521_o = n3504_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3523_o = n3504_o ? n3516_o : 1'b1;
  assign n3524_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3525_o = n3504_o ? 1'b1 : n3524_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3527_o = n3491_o ? 2'b01 : n3518_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3529_o = n3491_o ? 1'b0 : n3521_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3530_o = n3491_o ? n3503_o : n3523_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3531_o = n3491_o ? 1'b1 : n3525_o;
  /* TG68KdotC_Kernel.vhd:2027:66  */
  assign n3532_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2027:80  */
  assign n3533_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2027:74  */
  assign n3534_o = n3532_o | n3533_o;
  /* TG68KdotC_Kernel.vhd:2028:91  */
  assign n3535_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2028:103  */
  assign n3537_o = n3535_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2028:82  */
  assign n3538_o = nextpass | n3537_o;
  /* TG68KdotC_Kernel.vhd:2028:118  */
  assign n3539_o = exec[31];
  /* TG68KdotC_Kernel.vhd:2028:126  */
  assign n3540_o = ~n3539_o;
  /* TG68KdotC_Kernel.vhd:2028:110  */
  assign n3541_o = n3540_o & n3538_o;
  /* TG68KdotC_Kernel.vhd:2028:146  */
  assign n3543_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2028:131  */
  assign n3544_o = n3543_o & n3541_o;
  /* TG68KdotC_Kernel.vhd:2028:65  */
  assign n3547_o = n3544_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:65  */
  assign n3551_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:65  */
  assign n3554_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3556_o = n3534_o ? n3551_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3558_o = n3534_o ? n3554_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3561_o = n3534_o ? 1'b1 : 1'b0;
  assign n3562_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3563_o = n3580_o ? 1'b1 : n3562_o;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3565_o = n3534_o ? n3547_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3566_o = n3490_o ? n3527_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3568_o = n3490_o ? n3556_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3570_o = n3490_o ? n3558_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3572_o = n3490_o ? n3529_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3574_o = n3490_o ? n3530_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3576_o = n3490_o ? n3561_o : 1'b0;
  assign n3577_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3578_o = n3490_o ? n3531_o : n3577_o;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3580_o = n3534_o & n3490_o;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3582_o = n3490_o ? n3565_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3583_o = n3357_o ? n1921_o : n3566_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3584_o = n3357_o ? n3457_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3586_o = n3357_o ? n3459_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3588_o = n3357_o ? n3461_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3589_o = n3357_o ? n3462_o : n3568_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3591_o = n3357_o ? n3464_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3592_o = n3357_o ? n3466_o : n3570_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3593_o = n3357_o ? n3467_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3594_o = n3357_o ? n3468_o : n3572_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3595_o = n3357_o ? n3469_o : n3574_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3596_o = n3357_o ? n3471_o : n3576_o;
  assign n3597_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3598_o = n3357_o ? n3597_o : n3578_o;
  assign n3599_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3600_o = n3357_o ? n3473_o : n3599_o;
  assign n3601_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3602_o = n3357_o ? n3601_o : n3563_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3604_o = n3357_o ? n3474_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3606_o = n3357_o ? n3476_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3608_o = n3357_o ? 1'b0 : n3582_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3610_o = n3357_o ? n3477_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3612_o = n3357_o ? n3479_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2044:52  */
  assign n3613_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:2046:67  */
  assign n3614_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2046:79  */
  assign n3616_o = n3614_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2047:67  */
  assign n3617_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2047:79  */
  assign n3619_o = n3617_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2047:96  */
  assign n3620_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2047:108  */
  assign n3622_o = n3620_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2047:87  */
  assign n3623_o = n3619_o | n3622_o;
  /* TG68KdotC_Kernel.vhd:2046:87  */
  assign n3624_o = n3623_o & n3616_o;
  /* TG68KdotC_Kernel.vhd:2048:74  */
  assign n3625_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2048:86  */
  assign n3627_o = n3625_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2049:93  */
  assign n3628_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2049:96  */
  assign n3629_o = ~n3628_o;
  /* TG68KdotC_Kernel.vhd:2049:101  */
  assign n3631_o = 1'b1 & n3629_o;
  /* TG68KdotC_Kernel.vhd:2049:86  */
  assign n3633_o = 1'b0 | n3631_o;
  /* TG68KdotC_Kernel.vhd:2049:116  */
  assign n3634_o = n3633_o | svmode;
  /* TG68KdotC_Kernel.vhd:2054:87  */
  assign n3636_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2054:104  */
  assign n3638_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2054:95  */
  assign n3639_o = n3638_o & n3636_o;
  /* TG68KdotC_Kernel.vhd:2054:123  */
  assign n3640_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2054:110  */
  assign n3641_o = n3640_o & n3639_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3643_o = n3705_o ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2057:90  */
  assign n3644_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2057:102  */
  assign n3646_o = n3644_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2057:81  */
  assign n3649_o = n3646_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2049:73  */
  assign n3650_o = n3641_o & n3634_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3652_o = n3706_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2049:73  */
  assign n3655_o = n3634_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2049:73  */
  assign n3658_o = n3634_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2049:73  */
  assign n3661_o = n3634_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2049:73  */
  assign n3664_o = n3634_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2049:73  */
  assign n3666_o = n3634_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2049:73  */
  assign n3668_o = n3634_o ? n3649_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2071:82  */
  assign n3672_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2071:94  */
  assign n3674_o = n3672_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2071:73  */
  assign n3677_o = n3674_o ? 1'b1 : 1'b0;
  assign n3679_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2074:73  */
  assign n3680_o = setexecopc ? 1'b1 : n3679_o;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3681_o = n3650_o & n3627_o;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3682_o = n3634_o & n3627_o;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3684_o = n3627_o ? n3655_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3687_o = n3627_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3689_o = n3627_o ? n3658_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3691_o = n3627_o ? n3661_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3693_o = n3627_o ? n3664_o : 1'b1;
  assign n3694_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3695_o = n3627_o ? n3694_o : n3680_o;
  assign n3696_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3697_o = n3627_o ? n3696_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3699_o = n3627_o ? n3666_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3701_o = n3627_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3703_o = n3627_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3704_o = n3627_o ? n3668_o : n3677_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3705_o = n3681_o & n3624_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3706_o = n3682_o & n3624_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3708_o = n3624_o ? n3684_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3710_o = n3624_o ? n3687_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3713_o = n3624_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3715_o = n3624_o ? n3689_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3717_o = n3624_o ? n3691_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3719_o = n3624_o ? n3693_o : 1'b0;
  assign n3720_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3721_o = n3624_o ? n3695_o : n3720_o;
  assign n3722_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3723_o = n3624_o ? n3697_o : n3722_o;
  assign n3724_o = {n3701_o, n3699_o};
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3726_o = n3624_o ? n3724_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3728_o = n3624_o ? n3703_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3730_o = n3624_o ? n3704_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2045:49  */
  assign n3732_o = n3613_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2083:67  */
  assign n3733_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2083:79  */
  assign n3735_o = n3733_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2084:67  */
  assign n3736_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2084:79  */
  assign n3738_o = n3736_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2084:96  */
  assign n3739_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2084:108  */
  assign n3741_o = n3739_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2084:87  */
  assign n3742_o = n3738_o | n3741_o;
  /* TG68KdotC_Kernel.vhd:2083:87  */
  assign n3743_o = n3742_o & n3735_o;
  /* TG68KdotC_Kernel.vhd:2085:74  */
  assign n3744_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2085:86  */
  assign n3746_o = n3744_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2086:93  */
  assign n3747_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2086:101  */
  assign n3749_o = 1'b1 & n3747_o;
  /* TG68KdotC_Kernel.vhd:2086:86  */
  assign n3751_o = 1'b0 | n3749_o;
  /* TG68KdotC_Kernel.vhd:2094:90  */
  assign n3753_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2094:102  */
  assign n3755_o = n3753_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2094:81  */
  assign n3758_o = n3755_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3760_o = n3813_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2086:73  */
  assign n3763_o = n3751_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2086:73  */
  assign n3766_o = n3751_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2086:73  */
  assign n3769_o = n3751_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2086:73  */
  assign n3772_o = n3751_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2086:73  */
  assign n3774_o = n3751_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2086:73  */
  assign n3776_o = n3751_o ? n3758_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2105:71  */
  assign n3778_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2105:88  */
  assign n3780_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2105:79  */
  assign n3781_o = n3780_o & n3778_o;
  /* TG68KdotC_Kernel.vhd:2105:107  */
  assign n3782_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2105:94  */
  assign n3783_o = n3782_o & n3781_o;
  /* TG68KdotC_Kernel.vhd:2105:65  */
  assign n3785_o = n3783_o ? 1'b1 : make_berr;
  assign n3787_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2108:73  */
  assign n3788_o = setexecopc ? 1'b1 : n3787_o;
  /* TG68KdotC_Kernel.vhd:2111:82  */
  assign n3789_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2111:94  */
  assign n3791_o = n3789_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2111:73  */
  assign n3794_o = n3791_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3795_o = n3746_o ? make_berr : n3785_o;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3796_o = n3751_o & n3746_o;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3798_o = n3746_o ? n3763_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3800_o = n3746_o ? n3766_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3802_o = n3746_o ? n3769_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3804_o = n3746_o ? n3772_o : 1'b1;
  assign n3805_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3806_o = n3746_o ? n3805_o : n3788_o;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3808_o = n3746_o ? n3774_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3810_o = n3746_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3811_o = n3746_o ? n3776_o : n3794_o;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3812_o = n3743_o ? n3795_o : make_berr;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3813_o = n3796_o & n3743_o;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3815_o = n3743_o ? n3798_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3817_o = n3743_o ? n3800_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3819_o = n3743_o ? n3802_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3821_o = n3743_o ? n3804_o : 1'b0;
  assign n3822_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3823_o = n3743_o ? n3806_o : n3822_o;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3825_o = n3743_o ? n3808_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3827_o = n3743_o ? n3810_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3829_o = n3743_o ? n3811_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2082:49  */
  assign n3831_o = n3613_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2120:66  */
  assign n3832_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2120:78  */
  assign n3834_o = n3832_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2121:74  */
  assign n3835_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2121:86  */
  assign n3837_o = n3835_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2122:75  */
  assign n3838_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2122:87  */
  assign n3840_o = n3838_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2122:105  */
  assign n3841_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2122:117  */
  assign n3843_o = n3841_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2122:96  */
  assign n3844_o = n3840_o | n3843_o;
  /* TG68KdotC_Kernel.vhd:2121:94  */
  assign n3845_o = n3844_o & n3837_o;
  /* TG68KdotC_Kernel.vhd:2126:101  */
  assign n3846_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2126:113  */
  assign n3848_o = n3846_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2126:91  */
  assign n3849_o = n3848_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2126:129  */
  assign n3851_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2126:148  */
  assign n3852_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2126:135  */
  assign n3853_o = n3852_o & n3851_o;
  /* TG68KdotC_Kernel.vhd:2126:120  */
  assign n3854_o = n3849_o | n3853_o;
  /* TG68KdotC_Kernel.vhd:2126:154  */
  assign n3855_o = n3854_o | direct_data;
  assign n3857_o = n1909_o[51];
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3858_o = n3928_o ? 1'b1 : n3857_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3860_o = n3920_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3863_o = n3845_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3866_o = n3845_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3869_o = n3845_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3872_o = n3845_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3874_o = n3855_o & n3845_o;
  /* TG68KdotC_Kernel.vhd:2134:75  */
  assign n3875_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2134:87  */
  assign n3877_o = n3875_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2135:75  */
  assign n3878_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2135:87  */
  assign n3880_o = n3878_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2135:104  */
  assign n3881_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2135:116  */
  assign n3883_o = n3881_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2135:95  */
  assign n3884_o = n3880_o | n3883_o;
  /* TG68KdotC_Kernel.vhd:2134:95  */
  assign n3885_o = n3884_o & n3877_o;
  /* TG68KdotC_Kernel.vhd:2141:82  */
  assign n3888_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2141:94  */
  assign n3890_o = n3888_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2141:73  */
  assign n3893_o = n3890_o ? 1'b1 : 1'b0;
  assign n3895_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3896_o = n3913_o ? 1'b1 : n3895_o;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3899_o = n3885_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3902_o = n3885_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3905_o = n3885_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3908_o = n3885_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3911_o = n3885_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3913_o = setexecopc & n3885_o;
  assign n3914_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3915_o = n3885_o ? 1'b1 : n3914_o;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3917_o = n3885_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3919_o = n3885_o ? n3893_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3920_o = n3845_o & n3834_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3922_o = n3834_o ? 1'b0 : n3899_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3923_o = n3834_o ? n3863_o : n3902_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3924_o = n3834_o ? n3866_o : n3905_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3925_o = n3834_o ? n3869_o : n3908_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3926_o = n3834_o ? n3872_o : n3911_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3928_o = n3874_o & n3834_o;
  assign n3929_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3930_o = n3834_o ? n3929_o : n3896_o;
  assign n3931_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3932_o = n3834_o ? n3931_o : n3915_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3934_o = n3834_o ? 1'b0 : n3917_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3936_o = n3834_o ? 1'b0 : n3919_o;
  /* TG68KdotC_Kernel.vhd:2119:49  */
  assign n3938_o = n3613_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:2153:66  */
  assign n3939_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2153:78  */
  assign n3941_o = n3939_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2154:74  */
  assign n3942_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2154:86  */
  assign n3944_o = n3942_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2155:75  */
  assign n3945_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2155:87  */
  assign n3947_o = n3945_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2155:105  */
  assign n3948_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2155:117  */
  assign n3950_o = n3948_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2155:96  */
  assign n3951_o = n3947_o | n3950_o;
  /* TG68KdotC_Kernel.vhd:2154:94  */
  assign n3952_o = n3951_o & n3944_o;
  /* TG68KdotC_Kernel.vhd:2160:109  */
  assign n3953_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2160:121  */
  assign n3955_o = n3953_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2160:99  */
  assign n3956_o = n3955_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2160:137  */
  assign n3958_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2160:156  */
  assign n3959_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2160:143  */
  assign n3960_o = n3959_o & n3958_o;
  /* TG68KdotC_Kernel.vhd:2160:128  */
  assign n3961_o = n3956_o | n3960_o;
  /* TG68KdotC_Kernel.vhd:2160:162  */
  assign n3962_o = n3961_o | direct_data;
  assign n3965_o = {1'b1, 1'b1};
  assign n3966_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3967_o = n4068_o ? n3965_o : n3966_o;
  /* TG68KdotC_Kernel.vhd:2164:88  */
  assign n3968_o = exec[52];
  /* TG68KdotC_Kernel.vhd:2164:128  */
  assign n3969_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2164:140  */
  assign n3971_o = n3969_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2164:118  */
  assign n3972_o = n3971_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2164:100  */
  assign n3973_o = n3968_o | n3972_o;
  /* TG68KdotC_Kernel.vhd:2164:156  */
  assign n3975_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2164:175  */
  assign n3976_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2164:162  */
  assign n3977_o = n3976_o & n3975_o;
  /* TG68KdotC_Kernel.vhd:2164:147  */
  assign n3978_o = n3973_o | n3977_o;
  /* TG68KdotC_Kernel.vhd:2164:181  */
  assign n3979_o = n3978_o | direct_data;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3981_o = n4057_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3983_o = n4056_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3984_o = n3979_o & svmode;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3987_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3990_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3993_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3996_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3998_o = n3962_o & svmode;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3999_o = svmode & n3952_o;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n4000_o = n3984_o & n3952_o;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n4002_o = n3952_o ? n3987_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n4005_o = n3952_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n4007_o = n3952_o ? n3990_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n4009_o = n3952_o ? n3993_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n4011_o = n3952_o ? n3996_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n4013_o = n3998_o & n3952_o;
  /* TG68KdotC_Kernel.vhd:2176:74  */
  assign n4014_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2176:86  */
  assign n4016_o = n4014_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2177:75  */
  assign n4017_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2177:87  */
  assign n4019_o = n4017_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2177:104  */
  assign n4020_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2177:116  */
  assign n4022_o = n4020_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2177:95  */
  assign n4023_o = n4019_o | n4022_o;
  /* TG68KdotC_Kernel.vhd:2176:94  */
  assign n4024_o = n4023_o & n4016_o;
  /* TG68KdotC_Kernel.vhd:2182:82  */
  assign n4027_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2182:94  */
  assign n4029_o = n4027_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2182:73  */
  assign n4032_o = n4029_o ? 1'b1 : 1'b0;
  assign n4034_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4035_o = n4049_o ? 1'b1 : n4034_o;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4038_o = n4024_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4041_o = n4024_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4044_o = n4024_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4047_o = n4024_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4049_o = setexecopc & n4024_o;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4051_o = n4024_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4053_o = n4024_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n4055_o = n4024_o ? n4032_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4056_o = n3999_o & n3941_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4057_o = n4000_o & n3941_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4059_o = n3941_o ? 1'b0 : n4038_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4061_o = n3941_o ? n4002_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4062_o = n3941_o ? n4005_o : n4041_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4064_o = n3941_o ? n4007_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4065_o = n3941_o ? n4009_o : n4044_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4066_o = n3941_o ? n4011_o : n4047_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4068_o = n4013_o & n3941_o;
  assign n4069_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4070_o = n3941_o ? n4069_o : n4035_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4072_o = n3941_o ? 1'b0 : n4051_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4074_o = n3941_o ? 1'b0 : n4053_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4076_o = n3941_o ? 1'b0 : n4055_o;
  /* TG68KdotC_Kernel.vhd:2152:49  */
  assign n4078_o = n3613_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:2194:66  */
  assign n4079_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2195:74  */
  assign n4080_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2195:86  */
  assign n4082_o = n4080_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2195:103  */
  assign n4083_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2195:107  */
  assign n4084_o = ~n4083_o;
  /* TG68KdotC_Kernel.vhd:2195:93  */
  assign n4085_o = n4084_o & n4082_o;
  /* TG68KdotC_Kernel.vhd:2200:82  */
  assign n4089_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2200:85  */
  assign n4090_o = ~n4089_o;
  /* TG68KdotC_Kernel.vhd:2200:73  */
  assign n4093_o = n4090_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2200:73  */
  assign n4095_o = n4090_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:83  */
  assign n4096_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2206:103  */
  assign n4097_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:2206:120  */
  assign n4098_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:2206:132  */
  assign n4100_o = n4098_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2206:111  */
  assign n4101_o = n4097_o | n4100_o;
  /* TG68KdotC_Kernel.vhd:2207:83  */
  assign n4102_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2207:95  */
  assign n4104_o = n4102_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2207:112  */
  assign n4105_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2207:124  */
  assign n4107_o = n4105_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2207:103  */
  assign n4108_o = n4104_o | n4107_o;
  /* TG68KdotC_Kernel.vhd:2206:139  */
  assign n4109_o = n4108_o & n4101_o;
  /* TG68KdotC_Kernel.vhd:2206:92  */
  assign n4110_o = n4096_o | n4109_o;
  /* TG68KdotC_Kernel.vhd:2208:83  */
  assign n4111_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2208:87  */
  assign n4112_o = ~n4111_o;
  /* TG68KdotC_Kernel.vhd:2208:102  */
  assign n4113_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2208:114  */
  assign n4115_o = n4113_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2209:82  */
  assign n4116_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2209:94  */
  assign n4118_o = n4116_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:2208:121  */
  assign n4119_o = n4118_o & n4115_o;
  /* TG68KdotC_Kernel.vhd:2210:82  */
  assign n4120_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2210:94  */
  assign n4122_o = n4120_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2209:102  */
  assign n4123_o = n4122_o & n4119_o;
  /* TG68KdotC_Kernel.vhd:2208:92  */
  assign n4124_o = n4112_o | n4123_o;
  /* TG68KdotC_Kernel.vhd:2207:133  */
  assign n4125_o = n4124_o & n4110_o;
  /* TG68KdotC_Kernel.vhd:2213:90  */
  assign n4127_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2213:93  */
  assign n4128_o = ~n4127_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4130_o = n4218_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2216:91  */
  assign n4131_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2216:103  */
  assign n4133_o = n4131_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2216:119  */
  assign n4134_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2216:131  */
  assign n4136_o = n4134_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:2216:110  */
  assign n4137_o = n4133_o | n4136_o;
  /* TG68KdotC_Kernel.vhd:2216:148  */
  assign n4139_o = state == 2'b01;
  /* TG68KdotC_Kernel.vhd:2216:139  */
  assign n4140_o = n4139_o & n4137_o;
  /* TG68KdotC_Kernel.vhd:2216:81  */
  assign n4144_o = n4140_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2216:81  */
  assign n4146_o = n4140_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2220:90  */
  assign n4147_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2220:102  */
  assign n4149_o = n4147_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2220:81  */
  assign n4153_o = n4149_o ? 1'b1 : 1'b0;
  assign n4154_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:2220:81  */
  assign n4155_o = n4149_o ? 1'b1 : n4154_o;
  /* TG68KdotC_Kernel.vhd:2224:89  */
  assign n4157_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2224:108  */
  assign n4158_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2224:95  */
  assign n4159_o = n4158_o & n4157_o;
  assign n4162_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4163_o = n4233_o ? 1'b1 : n4162_o;
  assign n4164_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4165_o = n4235_o ? 1'b1 : n4164_o;
  /* TG68KdotC_Kernel.vhd:2230:98  */
  assign n4167_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2230:110  */
  assign n4169_o = n4167_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:2230:126  */
  assign n4170_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2230:138  */
  assign n4172_o = n4170_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:2230:117  */
  assign n4173_o = n4169_o | n4172_o;
  /* TG68KdotC_Kernel.vhd:2230:154  */
  assign n4174_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2230:166  */
  assign n4176_o = n4174_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2230:145  */
  assign n4177_o = n4173_o | n4176_o;
  assign n4179_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2230:89  */
  assign n4180_o = n4177_o ? n4179_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2230:89  */
  assign n4183_o = n4177_o ? 7'b0011010 : 7'b0000001;
  assign n4184_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4185_o = n4239_o ? n4180_o : n4184_o;
  assign n4186_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4187_o = n4246_o ? 1'b1 : n4186_o;
  /* TG68KdotC_Kernel.vhd:2228:81  */
  assign n4188_o = decodeopc ? n4183_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2237:87  */
  assign n4189_o = set[62];
  /* TG68KdotC_Kernel.vhd:2240:106  */
  assign n4191_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2240:110  */
  assign n4192_o = ~n4191_o;
  /* TG68KdotC_Kernel.vhd:2240:97  */
  assign n4196_o = n4192_o ? 2'b11 : 2'b10;
  assign n4197_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4198_o = n4237_o ? 1'b1 : n4197_o;
  /* TG68KdotC_Kernel.vhd:2238:89  */
  assign n4201_o = movem_run ? n4196_o : 2'b01;
  /* TG68KdotC_Kernel.vhd:2238:89  */
  assign n4203_o = n4192_o & movem_run;
  assign n4204_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4205_o = n4242_o ? 1'b1 : n4204_o;
  assign n4206_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4207_o = n4244_o ? 1'b1 : n4206_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4209_o = n4217_o ? 7'b0011011 : n4188_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4210_o = n4219_o ? n4201_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4212_o = n4203_o & n4189_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4214_o = movem_run & n4189_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4216_o = movem_run & n4189_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4217_o = movem_run & n4189_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4218_o = n4128_o & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4219_o = n4189_o & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4222_o = n4125_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4224_o = n4125_o ? n4153_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4227_o = n4125_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4230_o = n4125_o ? 1'b0 : 1'b1;
  assign n4231_o = {1'b1, n4155_o};
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4233_o = n4159_o & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4235_o = n4159_o & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4237_o = n4212_o & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4239_o = decodeopc & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4240_o = n4125_o ? n4231_o : n2177_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4242_o = n4214_o & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4244_o = n4216_o & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4246_o = decodeopc & n4125_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4248_o = n4125_o ? n4144_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4250_o = n4125_o ? n4146_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4251_o = n4125_o ? n4209_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4252_o = n4085_o ? n4093_o : n4130_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4253_o = n4085_o ? n2026_o : n4210_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4255_o = n4085_o ? 1'b0 : n4222_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4258_o = n4085_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4260_o = n4085_o ? 1'b0 : n4224_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4262_o = n4085_o ? 1'b0 : n4227_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4264_o = n4085_o ? 1'b0 : n4230_o;
  assign n4265_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4266_o = n4085_o ? n4265_o : n4163_o;
  assign n4267_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4268_o = n4085_o ? n4267_o : n4165_o;
  assign n4269_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4270_o = n4085_o ? n4269_o : n4198_o;
  assign n4271_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4272_o = n4085_o ? n4271_o : n4185_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4273_o = n4085_o ? n2177_o : n4240_o;
  assign n4274_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4275_o = n4085_o ? n4274_o : n4205_o;
  assign n4276_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4277_o = n4085_o ? n4276_o : n4207_o;
  assign n4278_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4279_o = n4085_o ? n4278_o : n4187_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4281_o = n4085_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4283_o = n4085_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4285_o = n4085_o ? 1'b0 : n4248_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4286_o = n4085_o ? 1'b1 : n4250_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4288_o = n4085_o ? n4095_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4289_o = n4085_o ? n2180_o : n4251_o;
  /* TG68KdotC_Kernel.vhd:2258:74  */
  assign n4290_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2260:82  */
  assign n4291_o = opcode[8:7];
  /* TG68KdotC_Kernel.vhd:2260:94  */
  assign n4293_o = n4291_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2260:110  */
  assign n4294_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2260:122  */
  assign n4296_o = n4294_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2260:100  */
  assign n4297_o = n4296_o & n4293_o;
  /* TG68KdotC_Kernel.vhd:2260:141  */
  assign n4298_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2260:153  */
  assign n4300_o = n4298_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2260:171  */
  assign n4301_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2260:183  */
  assign n4303_o = n4301_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2260:162  */
  assign n4304_o = n4300_o | n4303_o;
  /* TG68KdotC_Kernel.vhd:2260:130  */
  assign n4305_o = n4304_o & n4297_o;
  /* TG68KdotC_Kernel.vhd:2260:190  */
  assign n4307_o = 1'b1 & n4305_o;
  /* TG68KdotC_Kernel.vhd:2261:102  */
  assign n4308_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2261:105  */
  assign n4309_o = ~n4308_o;
  /* TG68KdotC_Kernel.vhd:2261:133  */
  assign n4310_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2261:141  */
  assign n4312_o = 1'b1 & n4310_o;
  /* TG68KdotC_Kernel.vhd:2261:126  */
  assign n4314_o = 1'b0 | n4312_o;
  /* TG68KdotC_Kernel.vhd:2261:110  */
  assign n4315_o = n4314_o & n4309_o;
  /* TG68KdotC_Kernel.vhd:2261:91  */
  assign n4316_o = n4315_o & n4307_o;
  assign n4319_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2262:81  */
  assign n4320_o = decodeopc ? 1'b1 : n4319_o;
  assign n4321_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2262:81  */
  assign n4322_o = decodeopc ? 1'b1 : n4321_o;
  /* TG68KdotC_Kernel.vhd:2262:81  */
  assign n4324_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2267:96  */
  assign n4326_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2267:102  */
  assign n4327_o = nextpass & n4326_o;
  /* TG68KdotC_Kernel.vhd:2267:130  */
  assign n4328_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2267:142  */
  assign n4330_o = n4328_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2267:156  */
  assign n4331_o = exec[42];
  /* TG68KdotC_Kernel.vhd:2267:148  */
  assign n4332_o = n4331_o & n4330_o;
  /* TG68KdotC_Kernel.vhd:2267:120  */
  assign n4333_o = n4327_o | n4332_o;
  /* TG68KdotC_Kernel.vhd:2272:98  */
  assign n4336_o = sndopc[10];
  /* TG68KdotC_Kernel.vhd:2267:81  */
  assign n4338_o = n4344_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2267:81  */
  assign n4340_o = n4354_o ? 7'b1010100 : n4324_o;
  /* TG68KdotC_Kernel.vhd:2267:81  */
  assign n4344_o = n4336_o & n4333_o;
  /* TG68KdotC_Kernel.vhd:2267:81  */
  assign n4347_o = n4333_o ? 1'b1 : 1'b0;
  assign n4348_o = n1909_o[20];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4349_o = n4750_o ? 1'b1 : n4348_o;
  assign n4350_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4351_o = n4754_o ? 1'b1 : n4350_o;
  assign n4352_o = n1909_o[67];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4353_o = n4770_o ? 1'b1 : n4352_o;
  /* TG68KdotC_Kernel.vhd:2267:81  */
  assign n4354_o = n4336_o & n4333_o;
  /* TG68KdotC_Kernel.vhd:2282:85  */
  assign n4355_o = opcode[8:7];
  /* TG68KdotC_Kernel.vhd:2282:97  */
  assign n4357_o = n4355_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2282:113  */
  assign n4358_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2282:125  */
  assign n4360_o = n4358_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2282:103  */
  assign n4361_o = n4360_o & n4357_o;
  /* TG68KdotC_Kernel.vhd:2282:144  */
  assign n4362_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2282:156  */
  assign n4364_o = n4362_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2282:174  */
  assign n4365_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2282:186  */
  assign n4367_o = n4365_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2282:165  */
  assign n4368_o = n4364_o | n4367_o;
  /* TG68KdotC_Kernel.vhd:2282:133  */
  assign n4369_o = n4368_o & n4361_o;
  /* TG68KdotC_Kernel.vhd:2283:84  */
  assign n4370_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2283:115  */
  assign n4371_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2283:123  */
  assign n4373_o = 1'b1 & n4371_o;
  /* TG68KdotC_Kernel.vhd:2283:108  */
  assign n4375_o = 1'b0 | n4373_o;
  /* TG68KdotC_Kernel.vhd:2283:92  */
  assign n4376_o = n4375_o & n4370_o;
  /* TG68KdotC_Kernel.vhd:2284:83  */
  assign n4377_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2284:86  */
  assign n4378_o = ~n4377_o;
  /* TG68KdotC_Kernel.vhd:2284:114  */
  assign n4379_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2284:122  */
  assign n4381_o = 1'b1 & n4379_o;
  /* TG68KdotC_Kernel.vhd:2284:107  */
  assign n4383_o = 1'b0 | n4381_o;
  /* TG68KdotC_Kernel.vhd:2284:91  */
  assign n4384_o = n4383_o & n4378_o;
  /* TG68KdotC_Kernel.vhd:2283:141  */
  assign n4385_o = n4376_o | n4384_o;
  /* TG68KdotC_Kernel.vhd:2282:193  */
  assign n4386_o = n4385_o & n4369_o;
  assign n4389_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4390_o = n4451_o ? 1'b1 : n4389_o;
  assign n4391_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4392_o = n4453_o ? 1'b1 : n4391_o;
  /* TG68KdotC_Kernel.vhd:2285:81  */
  assign n4394_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2290:96  */
  assign n4396_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2290:102  */
  assign n4397_o = nextpass & n4396_o;
  /* TG68KdotC_Kernel.vhd:2290:130  */
  assign n4398_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2290:142  */
  assign n4400_o = n4398_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2290:156  */
  assign n4401_o = exec[42];
  /* TG68KdotC_Kernel.vhd:2290:148  */
  assign n4402_o = n4401_o & n4400_o;
  /* TG68KdotC_Kernel.vhd:2290:120  */
  assign n4403_o = n4397_o | n4402_o;
  /* TG68KdotC_Kernel.vhd:2294:98  */
  assign n4404_o = opcode[6];
  assign n4406_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2294:89  */
  assign n4407_o = n4404_o ? n4406_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2294:89  */
  assign n4410_o = n4404_o ? 7'b1010101 : 7'b1010001;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4412_o = n4432_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2290:81  */
  assign n4415_o = n4403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2290:81  */
  assign n4418_o = n4403_o ? 1'b1 : 1'b0;
  assign n4419_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4420_o = n4449_o ? n4407_o : n4419_o;
  /* TG68KdotC_Kernel.vhd:2290:81  */
  assign n4421_o = n4403_o ? n4410_o : n4394_o;
  /* TG68KdotC_Kernel.vhd:2302:107  */
  assign n4422_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2302:119  */
  assign n4424_o = n4422_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2302:125  */
  assign n4425_o = decodeopc & n4424_o;
  /* TG68KdotC_Kernel.vhd:2302:97  */
  assign n4426_o = nextpass | n4425_o;
  /* TG68KdotC_Kernel.vhd:2302:81  */
  assign n4429_o = n4426_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4431_o = n4386_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4432_o = n4403_o & n4386_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4435_o = n4386_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4437_o = n4386_o ? n4415_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4439_o = n4386_o ? n4418_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4441_o = n4386_o ? n4429_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4444_o = n4386_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4447_o = n4386_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4449_o = n4403_o & n4386_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4451_o = decodeopc & n4386_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4453_o = decodeopc & n4386_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4454_o = n4386_o ? n4421_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4456_o = n4316_o ? 2'b10 : n4431_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4457_o = n4316_o ? n4338_o : n4412_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4459_o = n4316_o ? 1'b1 : n4435_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4461_o = n4316_o ? 1'b0 : n4437_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4462_o = n4316_o ? n4347_o : n4439_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4464_o = n4316_o ? 1'b0 : n4441_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4466_o = n4316_o ? 1'b0 : n4444_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4468_o = n4316_o ? 1'b0 : n4447_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4470_o = n4333_o & n4316_o;
  assign n4471_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4472_o = n4316_o ? n4471_o : n4420_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4474_o = n4333_o & n4316_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4475_o = n4316_o ? n4320_o : n4390_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4477_o = n4333_o & n4316_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4478_o = n4316_o ? n4322_o : n4392_o;
  /* TG68KdotC_Kernel.vhd:2260:73  */
  assign n4479_o = n4316_o ? n4340_o : n4454_o;
  /* TG68KdotC_Kernel.vhd:2312:82  */
  assign n4480_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2314:90  */
  assign n4481_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2314:102  */
  assign n4483_o = n4481_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2317:93  */
  assign n4486_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2317:105  */
  assign n4488_o = n4486_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2321:99  */
  assign n4489_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:2321:116  */
  assign n4490_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:2321:128  */
  assign n4492_o = n4490_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2321:107  */
  assign n4493_o = n4489_o | n4492_o;
  /* TG68KdotC_Kernel.vhd:2322:98  */
  assign n4494_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2322:110  */
  assign n4496_o = n4494_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:2321:135  */
  assign n4497_o = n4496_o & n4493_o;
  /* TG68KdotC_Kernel.vhd:2323:98  */
  assign n4498_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2323:110  */
  assign n4500_o = n4498_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2322:118  */
  assign n4501_o = n4500_o & n4497_o;
  /* TG68KdotC_Kernel.vhd:2326:128  */
  assign n4503_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2326:113  */
  assign n4504_o = n4503_o & nextpass;
  /* TG68KdotC_Kernel.vhd:2326:97  */
  assign n4507_o = n4504_o ? 2'b11 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4509_o = n4520_o ? 1'b1 : n2015_o;
  assign n4510_o = n2162_o[1];
  assign n4511_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4512_o = n2037_o ? n4510_o : n4511_o;
  /* TG68KdotC_Kernel.vhd:2326:97  */
  assign n4513_o = n4504_o ? 1'b1 : n4512_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4515_o = n4537_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2332:103  */
  assign n4516_o = set[62];
  /* TG68KdotC_Kernel.vhd:2332:97  */
  assign n4518_o = n4516_o ? 2'b01 : n4507_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4519_o = n4501_o ? n4518_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4520_o = n4504_o & n4501_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4523_o = n4501_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4526_o = n4501_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4529_o = n4501_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4532_o = n4501_o ? 1'b1 : 1'b0;
  assign n4533_o = n2162_o[1];
  assign n4534_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4535_o = n2037_o ? n4533_o : n4534_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4536_o = n4501_o ? n4513_o : n4535_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4537_o = n4504_o & n4501_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4538_o = n4488_o ? n2026_o : n4519_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4539_o = n4488_o ? n2015_o : n4509_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4541_o = n4488_o ? 1'b0 : n4523_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4543_o = n4488_o ? 1'b1 : n4526_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4545_o = n4488_o ? 1'b1 : n4529_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4547_o = n4488_o ? 1'b0 : n4532_o;
  assign n4548_o = n2162_o[1];
  assign n4549_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4550_o = n2037_o ? n4548_o : n4549_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4551_o = n4488_o ? n4550_o : n4536_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4552_o = n4488_o ? n2180_o : n4515_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4553_o = n4483_o ? n2026_o : n4538_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4554_o = n4483_o ? n2015_o : n4539_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4556_o = n4483_o ? 1'b0 : n4541_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4558_o = n4483_o ? 1'b0 : n4543_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4560_o = n4483_o ? 1'b0 : n4545_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4562_o = n4483_o ? 1'b0 : n4547_o;
  assign n4563_o = n2162_o[1];
  assign n4564_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4565_o = n2037_o ? n4563_o : n4564_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4566_o = n4483_o ? n4565_o : n4551_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4568_o = n4483_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4570_o = n4483_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4571_o = n4483_o ? n2180_o : n4552_o;
  /* TG68KdotC_Kernel.vhd:2341:90  */
  assign n4572_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2341:102  */
  assign n4574_o = n4572_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4584_o = n4659_o ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2346:89  */
  assign n4587_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2346:89  */
  assign n4590_o = decodeopc ? 1'b1 : 1'b0;
  assign n4591_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4592_o = n4670_o ? 1'b1 : n4591_o;
  assign n4593_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4594_o = n4672_o ? 1'b1 : n4593_o;
  assign n4595_o = n2162_o[1];
  assign n4596_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4597_o = n2037_o ? n4595_o : n4596_o;
  /* TG68KdotC_Kernel.vhd:2346:89  */
  assign n4598_o = decodeopc ? 1'b1 : n4597_o;
  assign n4599_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4600_o = n4682_o ? 1'b1 : n4599_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4601_o = n4685_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4603_o = n4692_o ? 7'b0100011 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2358:98  */
  assign n4604_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2358:110  */
  assign n4606_o = n4604_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2359:99  */
  assign n4607_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2359:111  */
  assign n4609_o = n4607_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2359:128  */
  assign n4610_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2359:140  */
  assign n4612_o = n4610_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2359:119  */
  assign n4613_o = n4609_o | n4612_o;
  /* TG68KdotC_Kernel.vhd:2358:118  */
  assign n4614_o = n4613_o & n4606_o;
  /* TG68KdotC_Kernel.vhd:2367:106  */
  assign n4619_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2367:118  */
  assign n4621_o = n4619_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2367:97  */
  assign n4624_o = n4621_o ? 1'b1 : 1'b0;
  assign n4626_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4627_o = n4644_o ? 1'b1 : n4626_o;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4630_o = n4614_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4633_o = n4614_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4636_o = n4614_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4639_o = n4614_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4642_o = n4614_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4644_o = setexecopc & n4614_o;
  assign n4645_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4646_o = n4614_o ? 1'b1 : n4645_o;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4648_o = n4614_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4650_o = n4614_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4652_o = n4614_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4654_o = n4614_o ? n4624_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4656_o = n4574_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4658_o = n4574_o ? 1'b0 : n4630_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4659_o = decodeopc & n4574_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4661_o = n4574_o ? n4587_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4662_o = n4574_o ? n4590_o : n4633_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4664_o = n4574_o ? 1'b0 : n4636_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4666_o = n4574_o ? 1'b0 : n4639_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4668_o = n4574_o ? 1'b0 : n4642_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4670_o = decodeopc & n4574_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4672_o = decodeopc & n4574_o;
  assign n4673_o = n2162_o[1];
  assign n4674_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4675_o = n2037_o ? n4673_o : n4674_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4676_o = n4574_o ? n4598_o : n4675_o;
  assign n4677_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4678_o = n4574_o ? 1'b1 : n4677_o;
  assign n4679_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4680_o = n4574_o ? n4679_o : n4627_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4682_o = decodeopc & n4574_o;
  assign n4683_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4684_o = n4574_o ? n4683_o : n4646_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4685_o = decodeopc & n4574_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4686_o = n4574_o ? 1'b1 : n4648_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4688_o = n4574_o ? 1'b0 : n4650_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4690_o = n4574_o ? 1'b0 : n4652_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4691_o = n4574_o ? 1'b1 : n4654_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4692_o = decodeopc & n4574_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4694_o = n4480_o ? 2'b10 : n4656_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4695_o = n4480_o ? n4553_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4697_o = n4480_o ? 1'b0 : n4658_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4698_o = n4480_o ? n4554_o : n4584_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4700_o = n4480_o ? n4556_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4702_o = n4480_o ? 1'b0 : n4661_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4704_o = n4480_o ? 1'b0 : n4662_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4705_o = n4480_o ? n4558_o : n4664_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4706_o = n4480_o ? n4560_o : n4666_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4707_o = n4480_o ? n4562_o : n4668_o;
  assign n4708_o = {n4684_o, n4600_o, n4680_o};
  assign n4709_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4710_o = n4480_o ? n4709_o : n4592_o;
  assign n4711_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4712_o = n4480_o ? n4711_o : n4594_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4713_o = n4480_o ? n4566_o : n4676_o;
  assign n4714_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4715_o = n4480_o ? n4714_o : n4678_o;
  assign n4716_o = n1909_o[56:54];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4717_o = n4480_o ? n4716_o : n4708_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4718_o = n4480_o ? n2171_o : n4601_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4720_o = n4480_o ? 1'b0 : n4686_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4722_o = n4480_o ? 1'b0 : n4688_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4724_o = n4480_o ? n4568_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4726_o = n4480_o ? 1'b0 : n4690_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4727_o = n4480_o ? n4570_o : n4691_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4728_o = n4480_o ? n4571_o : n4603_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4729_o = n4290_o ? n4456_o : n4694_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4730_o = n4290_o ? n4457_o : n4695_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4732_o = n4290_o ? 1'b0 : n4697_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4733_o = n4290_o ? n2015_o : n4698_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4735_o = n4290_o ? 1'b0 : n4700_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4737_o = n4290_o ? 1'b0 : n4702_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4738_o = n4290_o ? n4459_o : n4704_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4740_o = n4290_o ? n4461_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4742_o = n4290_o ? n4462_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4744_o = n4290_o ? n4464_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4745_o = n4290_o ? n4466_o : n4705_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4746_o = n4290_o ? n4468_o : n4706_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4748_o = n4290_o ? 1'b0 : n4707_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4750_o = n4470_o & n4290_o;
  assign n4751_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4752_o = n4290_o ? n4472_o : n4751_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4754_o = n4474_o & n4290_o;
  assign n4755_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4756_o = n4290_o ? n4755_o : n4710_o;
  assign n4757_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4758_o = n4290_o ? n4475_o : n4757_o;
  assign n4759_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4760_o = n4290_o ? n4759_o : n4712_o;
  assign n4761_o = n2162_o[1];
  assign n4762_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4763_o = n2037_o ? n4761_o : n4762_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4764_o = n4290_o ? n4763_o : n4713_o;
  assign n4765_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4766_o = n4290_o ? n4765_o : n4715_o;
  assign n4767_o = n1909_o[56:54];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4768_o = n4290_o ? n4767_o : n4717_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4770_o = n4477_o & n4290_o;
  assign n4771_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4772_o = n4290_o ? n4478_o : n4771_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4773_o = n4290_o ? n2171_o : n4718_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4775_o = n4290_o ? 1'b0 : n4720_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4777_o = n4290_o ? 1'b0 : n4722_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4779_o = n4290_o ? 1'b0 : n4724_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4781_o = n4290_o ? 1'b0 : n4726_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4783_o = n4290_o ? 1'b0 : n4727_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4784_o = n4290_o ? n4479_o : n4728_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4785_o = n4079_o ? n4252_o : n4729_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4786_o = n4079_o ? n4253_o : n4730_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4788_o = n4079_o ? 1'b0 : n4732_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4789_o = n4079_o ? n2015_o : n4733_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4790_o = n4079_o ? n4255_o : n4735_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4792_o = n4079_o ? 1'b0 : n4737_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4793_o = n4079_o ? n4258_o : n4738_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4795_o = n4079_o ? 1'b0 : n4740_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4797_o = n4079_o ? 1'b0 : n4742_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4799_o = n4079_o ? 1'b0 : n4744_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4801_o = n4079_o ? n4260_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4802_o = n4079_o ? n4262_o : n4745_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4803_o = n4079_o ? n4264_o : n4746_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4805_o = n4079_o ? 1'b0 : n4748_o;
  assign n4806_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4807_o = n4079_o ? n4266_o : n4806_o;
  assign n4808_o = n1909_o[20];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4809_o = n4079_o ? n4808_o : n4349_o;
  assign n4810_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4811_o = n4079_o ? n4810_o : n4752_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4812_o = n4079_o ? n4268_o : n4351_o;
  assign n4813_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4814_o = n4079_o ? n4813_o : n4756_o;
  assign n4815_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4816_o = n4079_o ? n4270_o : n4815_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4817_o = n4079_o ? n4272_o : n4758_o;
  assign n4818_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4819_o = n4079_o ? n4818_o : n4760_o;
  assign n4820_o = n2162_o[1];
  assign n4821_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4822_o = n2037_o ? n4820_o : n4821_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4823_o = n4079_o ? n4822_o : n4764_o;
  assign n4824_o = n4273_o[0];
  assign n4825_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4826_o = n4079_o ? n4824_o : n4825_o;
  assign n4827_o = n4273_o[1];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4828_o = n4079_o ? n4827_o : n4766_o;
  assign n4829_o = n4768_o[0];
  assign n4830_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4831_o = n4079_o ? n4830_o : n4829_o;
  assign n4832_o = n4768_o[1];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4833_o = n4079_o ? n4275_o : n4832_o;
  assign n4834_o = n4768_o[2];
  assign n4835_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4836_o = n4079_o ? n4835_o : n4834_o;
  assign n4837_o = n1909_o[67];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4838_o = n4079_o ? n4837_o : n4353_o;
  assign n4839_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4840_o = n4079_o ? n4277_o : n4839_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4841_o = n4079_o ? n4279_o : n4772_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4842_o = n4079_o ? n2171_o : n4773_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4844_o = n4079_o ? n4281_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4846_o = n4079_o ? 1'b0 : n4775_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4848_o = n4079_o ? n4283_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4850_o = n4079_o ? 1'b0 : n4777_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4852_o = n4079_o ? 1'b0 : n4779_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4854_o = n4079_o ? 1'b0 : n4781_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4856_o = n4079_o ? n4285_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4857_o = n4079_o ? n4286_o : n4783_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4859_o = n4079_o ? n4288_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4860_o = n4079_o ? n4289_o : n4784_o;
  /* TG68KdotC_Kernel.vhd:2193:49  */
  assign n4862_o = n3613_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2193:59  */
  assign n4864_o = n3613_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:2193:59  */
  assign n4865_o = n4862_o | n4864_o;
  /* TG68KdotC_Kernel.vhd:2384:66  */
  assign n4866_o = opcode[7:3];
  /* TG68KdotC_Kernel.vhd:2384:78  */
  assign n4868_o = n4866_o == 5'b11111;
  /* TG68KdotC_Kernel.vhd:2384:97  */
  assign n4869_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2384:109  */
  assign n4871_o = n4869_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2384:87  */
  assign n4872_o = n4871_o & n4868_o;
  /* TG68KdotC_Kernel.vhd:2388:75  */
  assign n4873_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2388:87  */
  assign n4875_o = n4873_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:2389:75  */
  assign n4876_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2389:87  */
  assign n4878_o = n4876_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2390:75  */
  assign n4879_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2390:87  */
  assign n4881_o = n4879_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2390:104  */
  assign n4882_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2390:116  */
  assign n4884_o = n4882_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2390:95  */
  assign n4885_o = n4881_o | n4884_o;
  /* TG68KdotC_Kernel.vhd:2389:95  */
  assign n4886_o = n4885_o & n4878_o;
  /* TG68KdotC_Kernel.vhd:2388:94  */
  assign n4887_o = n4875_o | n4886_o;
  /* TG68KdotC_Kernel.vhd:2391:76  */
  assign n4888_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2391:88  */
  assign n4890_o = n4888_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2391:105  */
  assign n4891_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2391:117  */
  assign n4893_o = n4891_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2391:95  */
  assign n4894_o = n4890_o | n4893_o;
  /* TG68KdotC_Kernel.vhd:2392:75  */
  assign n4895_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2392:87  */
  assign n4897_o = n4895_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2392:105  */
  assign n4898_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2392:117  */
  assign n4900_o = n4898_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2392:96  */
  assign n4901_o = n4897_o | n4900_o;
  /* TG68KdotC_Kernel.vhd:2391:127  */
  assign n4902_o = n4901_o & n4894_o;
  /* TG68KdotC_Kernel.vhd:2390:125  */
  assign n4903_o = n4902_o & n4887_o;
  /* TG68KdotC_Kernel.vhd:2396:90  */
  assign n4904_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2396:81  */
  assign n4907_o = n4904_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2394:73  */
  assign n4909_o = setexecopc ? n4907_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2394:73  */
  assign n4912_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2401:82  */
  assign n4914_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2401:94  */
  assign n4916_o = n4914_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2405:90  */
  assign n4917_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2405:102  */
  assign n4919_o = n4917_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2405:81  */
  assign n4922_o = n4919_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4924_o = n4933_o ? 2'b00 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2401:73  */
  assign n4927_o = n4916_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2401:73  */
  assign n4930_o = n4916_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2401:73  */
  assign n4932_o = n4916_o ? n4922_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4933_o = n4916_o & n4903_o;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4935_o = n4903_o ? n4927_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4937_o = n4903_o ? n4930_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4939_o = n4903_o ? n4909_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4941_o = n4903_o ? n4912_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4944_o = n4903_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4947_o = n4903_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4950_o = n4903_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4952_o = n4903_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4954_o = n4903_o ? n4932_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4955_o = n4872_o ? n1921_o : n4924_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4957_o = n4872_o ? 1'b0 : n4935_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4959_o = n4872_o ? 1'b0 : n4937_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4961_o = n4872_o ? 1'b0 : n4939_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4963_o = n4872_o ? 1'b0 : n4941_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4965_o = n4872_o ? 1'b1 : n4944_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4967_o = n4872_o ? 1'b1 : n4947_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4969_o = n4872_o ? 1'b0 : n4950_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4971_o = n4872_o ? 1'b0 : n4952_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4973_o = n4872_o ? 1'b0 : n4954_o;
  /* TG68KdotC_Kernel.vhd:2382:49  */
  assign n4975_o = n3613_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:2433:66  */
  assign n4976_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2434:75  */
  assign n4977_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:2434:92  */
  assign n4978_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:2434:104  */
  assign n4980_o = n4978_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2434:83  */
  assign n4981_o = n4977_o | n4980_o;
  /* TG68KdotC_Kernel.vhd:2435:74  */
  assign n4982_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2435:86  */
  assign n4984_o = n4982_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:2434:111  */
  assign n4985_o = n4984_o & n4981_o;
  /* TG68KdotC_Kernel.vhd:2435:104  */
  assign n4986_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2435:116  */
  assign n4988_o = n4986_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2435:94  */
  assign n4989_o = n4988_o & n4985_o;
  /* TG68KdotC_Kernel.vhd:2439:80  */
  assign n4990_o = exec[63];
  /* TG68KdotC_Kernel.vhd:2439:73  */
  assign n4992_o = n4990_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2442:104  */
  assign n4994_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2442:89  */
  assign n4995_o = n4994_o & nextpass;
  /* TG68KdotC_Kernel.vhd:2442:120  */
  assign n4996_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2442:123  */
  assign n4997_o = ~n4996_o;
  /* TG68KdotC_Kernel.vhd:2442:110  */
  assign n4998_o = n4997_o & n4995_o;
  /* TG68KdotC_Kernel.vhd:2442:73  */
  assign n5001_o = n4998_o ? 2'b11 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5003_o = n5039_o ? 1'b1 : n2015_o;
  assign n5004_o = n2162_o[1];
  assign n5005_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5006_o = n2037_o ? n5004_o : n5005_o;
  /* TG68KdotC_Kernel.vhd:2442:73  */
  assign n5007_o = n4998_o ? 1'b1 : n5006_o;
  /* TG68KdotC_Kernel.vhd:2442:73  */
  assign n5009_o = n4998_o ? 7'b0011000 : n4992_o;
  /* TG68KdotC_Kernel.vhd:2449:87  */
  assign n5011_o = micro_state == 7'b0000101;
  /* TG68KdotC_Kernel.vhd:2449:106  */
  assign n5012_o = brief[8];
  /* TG68KdotC_Kernel.vhd:2449:109  */
  assign n5013_o = ~n5012_o;
  /* TG68KdotC_Kernel.vhd:2449:97  */
  assign n5014_o = n5013_o & n5011_o;
  /* TG68KdotC_Kernel.vhd:2449:73  */
  assign n5016_o = n5014_o ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2452:81  */
  assign n5018_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:2452:73  */
  assign n5021_o = n5018_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2456:79  */
  assign n5023_o = set[62];
  /* TG68KdotC_Kernel.vhd:2457:88  */
  assign n5024_o = exec[73];
  /* TG68KdotC_Kernel.vhd:2457:100  */
  assign n5025_o = ~n5024_o;
  /* TG68KdotC_Kernel.vhd:2457:105  */
  assign n5026_o = n5025_o | long_done;
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n5028_o = n5030_o ? 1'b1 : n5016_o;
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n5030_o = n5026_o & n5023_o;
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n5032_o = n5023_o ? 2'b01 : n5001_o;
  assign n5033_o = n1909_o[63];
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n5034_o = n5023_o ? 1'b1 : n5033_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5035_o = n4989_o ? n5028_o : make_berr;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5037_o = n4989_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5038_o = n4989_o ? n5032_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5039_o = n4998_o & n4989_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5041_o = n4989_o ? n5021_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5044_o = n4989_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5047_o = n4989_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5050_o = n4989_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5053_o = n4989_o ? 1'b1 : 1'b0;
  assign n5054_o = {1'b1, n5034_o};
  assign n5055_o = n2162_o[1];
  assign n5056_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5057_o = n2037_o ? n5055_o : n5056_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5058_o = n4989_o ? n5007_o : n5057_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5059_o = n5607_o ? n5054_o : n2178_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n5060_o = n4989_o ? n5009_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2468:76  */
  assign n5061_o = opcode[6:0];
  /* TG68KdotC_Kernel.vhd:2469:73  */
  assign n5063_o = n5061_o == 7'b1000000;
  /* TG68KdotC_Kernel.vhd:2469:87  */
  assign n5065_o = n5061_o == 7'b1000001;
  /* TG68KdotC_Kernel.vhd:2469:87  */
  assign n5066_o = n5063_o | n5065_o;
  /* TG68KdotC_Kernel.vhd:2469:97  */
  assign n5068_o = n5061_o == 7'b1000010;
  /* TG68KdotC_Kernel.vhd:2469:97  */
  assign n5069_o = n5066_o | n5068_o;
  /* TG68KdotC_Kernel.vhd:2469:107  */
  assign n5071_o = n5061_o == 7'b1000011;
  /* TG68KdotC_Kernel.vhd:2469:107  */
  assign n5072_o = n5069_o | n5071_o;
  /* TG68KdotC_Kernel.vhd:2469:117  */
  assign n5074_o = n5061_o == 7'b1000100;
  /* TG68KdotC_Kernel.vhd:2469:117  */
  assign n5075_o = n5072_o | n5074_o;
  /* TG68KdotC_Kernel.vhd:2469:127  */
  assign n5077_o = n5061_o == 7'b1000101;
  /* TG68KdotC_Kernel.vhd:2469:127  */
  assign n5078_o = n5075_o | n5077_o;
  /* TG68KdotC_Kernel.vhd:2469:137  */
  assign n5080_o = n5061_o == 7'b1000110;
  /* TG68KdotC_Kernel.vhd:2469:137  */
  assign n5081_o = n5078_o | n5080_o;
  /* TG68KdotC_Kernel.vhd:2469:147  */
  assign n5083_o = n5061_o == 7'b1000111;
  /* TG68KdotC_Kernel.vhd:2469:147  */
  assign n5084_o = n5081_o | n5083_o;
  /* TG68KdotC_Kernel.vhd:2469:157  */
  assign n5086_o = n5061_o == 7'b1001000;
  /* TG68KdotC_Kernel.vhd:2469:157  */
  assign n5087_o = n5084_o | n5086_o;
  /* TG68KdotC_Kernel.vhd:2470:87  */
  assign n5089_o = n5061_o == 7'b1001001;
  /* TG68KdotC_Kernel.vhd:2470:87  */
  assign n5090_o = n5087_o | n5089_o;
  /* TG68KdotC_Kernel.vhd:2470:97  */
  assign n5092_o = n5061_o == 7'b1001010;
  /* TG68KdotC_Kernel.vhd:2470:97  */
  assign n5093_o = n5090_o | n5092_o;
  /* TG68KdotC_Kernel.vhd:2470:107  */
  assign n5095_o = n5061_o == 7'b1001011;
  /* TG68KdotC_Kernel.vhd:2470:107  */
  assign n5096_o = n5093_o | n5095_o;
  /* TG68KdotC_Kernel.vhd:2470:117  */
  assign n5098_o = n5061_o == 7'b1001100;
  /* TG68KdotC_Kernel.vhd:2470:117  */
  assign n5099_o = n5096_o | n5098_o;
  /* TG68KdotC_Kernel.vhd:2470:127  */
  assign n5101_o = n5061_o == 7'b1001101;
  /* TG68KdotC_Kernel.vhd:2470:127  */
  assign n5102_o = n5099_o | n5101_o;
  /* TG68KdotC_Kernel.vhd:2470:137  */
  assign n5104_o = n5061_o == 7'b1001110;
  /* TG68KdotC_Kernel.vhd:2470:137  */
  assign n5105_o = n5102_o | n5104_o;
  /* TG68KdotC_Kernel.vhd:2470:147  */
  assign n5107_o = n5061_o == 7'b1001111;
  /* TG68KdotC_Kernel.vhd:2470:147  */
  assign n5108_o = n5105_o | n5107_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n5116_o = decodeopc ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n5119_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n5122_o = decodeopc ? 1'b1 : 1'b0;
  assign n5123_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n5124_o = decodeopc ? 1'b1 : n5123_o;
  assign n5125_o = n2162_o[1];
  assign n5126_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5127_o = n2037_o ? n5125_o : n5126_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n5128_o = decodeopc ? 1'b1 : n5127_o;
  assign n5129_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n5130_o = decodeopc ? 1'b1 : n5129_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n5132_o = decodeopc ? 7'b0100011 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2474:73  */
  assign n5134_o = n5061_o == 7'b1010000;
  /* TG68KdotC_Kernel.vhd:2474:87  */
  assign n5136_o = n5061_o == 7'b1010001;
  /* TG68KdotC_Kernel.vhd:2474:87  */
  assign n5137_o = n5134_o | n5136_o;
  /* TG68KdotC_Kernel.vhd:2474:97  */
  assign n5139_o = n5061_o == 7'b1010010;
  /* TG68KdotC_Kernel.vhd:2474:97  */
  assign n5140_o = n5137_o | n5139_o;
  /* TG68KdotC_Kernel.vhd:2474:107  */
  assign n5142_o = n5061_o == 7'b1010011;
  /* TG68KdotC_Kernel.vhd:2474:107  */
  assign n5143_o = n5140_o | n5142_o;
  /* TG68KdotC_Kernel.vhd:2474:117  */
  assign n5145_o = n5061_o == 7'b1010100;
  /* TG68KdotC_Kernel.vhd:2474:117  */
  assign n5146_o = n5143_o | n5145_o;
  /* TG68KdotC_Kernel.vhd:2474:127  */
  assign n5148_o = n5061_o == 7'b1010101;
  /* TG68KdotC_Kernel.vhd:2474:127  */
  assign n5149_o = n5146_o | n5148_o;
  /* TG68KdotC_Kernel.vhd:2474:137  */
  assign n5151_o = n5061_o == 7'b1010110;
  /* TG68KdotC_Kernel.vhd:2474:137  */
  assign n5152_o = n5149_o | n5151_o;
  /* TG68KdotC_Kernel.vhd:2474:147  */
  assign n5154_o = n5061_o == 7'b1010111;
  /* TG68KdotC_Kernel.vhd:2474:147  */
  assign n5155_o = n5152_o | n5154_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5162_o = decodeopc ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5164_o = decodeopc ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5167_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5170_o = decodeopc ? 1'b1 : 1'b0;
  assign n5171_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5172_o = decodeopc ? 1'b1 : n5171_o;
  assign n5173_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5174_o = decodeopc ? 1'b1 : n5173_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5176_o = decodeopc ? 7'b0100101 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2489:73  */
  assign n5178_o = n5061_o == 7'b1011000;
  /* TG68KdotC_Kernel.vhd:2489:87  */
  assign n5180_o = n5061_o == 7'b1011001;
  /* TG68KdotC_Kernel.vhd:2489:87  */
  assign n5181_o = n5178_o | n5180_o;
  /* TG68KdotC_Kernel.vhd:2489:97  */
  assign n5183_o = n5061_o == 7'b1011010;
  /* TG68KdotC_Kernel.vhd:2489:97  */
  assign n5184_o = n5181_o | n5183_o;
  /* TG68KdotC_Kernel.vhd:2489:107  */
  assign n5186_o = n5061_o == 7'b1011011;
  /* TG68KdotC_Kernel.vhd:2489:107  */
  assign n5187_o = n5184_o | n5186_o;
  /* TG68KdotC_Kernel.vhd:2489:117  */
  assign n5189_o = n5061_o == 7'b1011100;
  /* TG68KdotC_Kernel.vhd:2489:117  */
  assign n5190_o = n5187_o | n5189_o;
  /* TG68KdotC_Kernel.vhd:2489:127  */
  assign n5192_o = n5061_o == 7'b1011101;
  /* TG68KdotC_Kernel.vhd:2489:127  */
  assign n5193_o = n5190_o | n5192_o;
  /* TG68KdotC_Kernel.vhd:2489:137  */
  assign n5195_o = n5061_o == 7'b1011110;
  /* TG68KdotC_Kernel.vhd:2489:137  */
  assign n5196_o = n5193_o | n5195_o;
  /* TG68KdotC_Kernel.vhd:2489:147  */
  assign n5198_o = n5061_o == 7'b1011111;
  /* TG68KdotC_Kernel.vhd:2489:147  */
  assign n5199_o = n5196_o | n5198_o;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5202_o = svmode ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5205_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5208_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5211_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5214_o = svmode ? 1'b0 : 1'b1;
  assign n5215_o = n2017_o[0];
  assign n5216_o = n1909_o[65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5217_o = n2010_o ? n5215_o : n5216_o;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5218_o = svmode ? 1'b1 : n5217_o;
  /* TG68KdotC_Kernel.vhd:2504:73  */
  assign n5220_o = n5061_o == 7'b1100000;
  /* TG68KdotC_Kernel.vhd:2504:87  */
  assign n5222_o = n5061_o == 7'b1100001;
  /* TG68KdotC_Kernel.vhd:2504:87  */
  assign n5223_o = n5220_o | n5222_o;
  /* TG68KdotC_Kernel.vhd:2504:97  */
  assign n5225_o = n5061_o == 7'b1100010;
  /* TG68KdotC_Kernel.vhd:2504:97  */
  assign n5226_o = n5223_o | n5225_o;
  /* TG68KdotC_Kernel.vhd:2504:107  */
  assign n5228_o = n5061_o == 7'b1100011;
  /* TG68KdotC_Kernel.vhd:2504:107  */
  assign n5229_o = n5226_o | n5228_o;
  /* TG68KdotC_Kernel.vhd:2504:117  */
  assign n5231_o = n5061_o == 7'b1100100;
  /* TG68KdotC_Kernel.vhd:2504:117  */
  assign n5232_o = n5229_o | n5231_o;
  /* TG68KdotC_Kernel.vhd:2504:127  */
  assign n5234_o = n5061_o == 7'b1100101;
  /* TG68KdotC_Kernel.vhd:2504:127  */
  assign n5235_o = n5232_o | n5234_o;
  /* TG68KdotC_Kernel.vhd:2504:137  */
  assign n5237_o = n5061_o == 7'b1100110;
  /* TG68KdotC_Kernel.vhd:2504:137  */
  assign n5238_o = n5235_o | n5237_o;
  /* TG68KdotC_Kernel.vhd:2504:147  */
  assign n5240_o = n5061_o == 7'b1100111;
  /* TG68KdotC_Kernel.vhd:2504:147  */
  assign n5241_o = n5238_o | n5240_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5245_o = svmode ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5248_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5251_o = svmode ? 1'b0 : 1'b1;
  assign n5252_o = n2017_o[1];
  assign n5253_o = n1909_o[66];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5254_o = n2010_o ? n5252_o : n5253_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5255_o = svmode ? 1'b1 : n5254_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5257_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2516:73  */
  assign n5259_o = n5061_o == 7'b1101000;
  /* TG68KdotC_Kernel.vhd:2516:87  */
  assign n5261_o = n5061_o == 7'b1101001;
  /* TG68KdotC_Kernel.vhd:2516:87  */
  assign n5262_o = n5259_o | n5261_o;
  /* TG68KdotC_Kernel.vhd:2516:97  */
  assign n5264_o = n5061_o == 7'b1101010;
  /* TG68KdotC_Kernel.vhd:2516:97  */
  assign n5265_o = n5262_o | n5264_o;
  /* TG68KdotC_Kernel.vhd:2516:107  */
  assign n5267_o = n5061_o == 7'b1101011;
  /* TG68KdotC_Kernel.vhd:2516:107  */
  assign n5268_o = n5265_o | n5267_o;
  /* TG68KdotC_Kernel.vhd:2516:117  */
  assign n5270_o = n5061_o == 7'b1101100;
  /* TG68KdotC_Kernel.vhd:2516:117  */
  assign n5271_o = n5268_o | n5270_o;
  /* TG68KdotC_Kernel.vhd:2516:127  */
  assign n5273_o = n5061_o == 7'b1101101;
  /* TG68KdotC_Kernel.vhd:2516:127  */
  assign n5274_o = n5271_o | n5273_o;
  /* TG68KdotC_Kernel.vhd:2516:137  */
  assign n5276_o = n5061_o == 7'b1101110;
  /* TG68KdotC_Kernel.vhd:2516:137  */
  assign n5277_o = n5274_o | n5276_o;
  /* TG68KdotC_Kernel.vhd:2516:147  */
  assign n5279_o = n5061_o == 7'b1101111;
  /* TG68KdotC_Kernel.vhd:2516:147  */
  assign n5280_o = n5277_o | n5279_o;
  /* TG68KdotC_Kernel.vhd:2528:90  */
  assign n5281_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:2533:89  */
  assign n5285_o = decodeopc ? 6'b000000 : n1906_o;
  assign n5286_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2533:89  */
  assign n5287_o = decodeopc ? 1'b1 : n5286_o;
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5288_o = n5281_o ? n1906_o : n5285_o;
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5291_o = n5281_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5294_o = n5281_o ? 1'b1 : 1'b0;
  assign n5295_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5296_o = n5281_o ? n5295_o : n5287_o;
  assign n5297_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5298_o = n5281_o ? n5297_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2527:73  */
  assign n5300_o = n5061_o == 7'b1110000;
  /* TG68KdotC_Kernel.vhd:2539:73  */
  assign n5302_o = n5061_o == 7'b1110001;
  /* TG68KdotC_Kernel.vhd:2542:90  */
  assign n5303_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:2546:89  */
  assign n5305_o = decodeopc ? 1'b1 : n2148_o;
  /* TG68KdotC_Kernel.vhd:2546:89  */
  assign n5308_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2550:89  */
  assign n5310_o = stop ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5311_o = n5303_o ? make_berr : n5310_o;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5312_o = n5303_o ? n2148_o : n5305_o;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5315_o = n5303_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5318_o = n5303_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5320_o = n5303_o ? 1'b0 : n5308_o;
  /* TG68KdotC_Kernel.vhd:2541:73  */
  assign n5322_o = n5061_o == 7'b1110010;
  /* TG68KdotC_Kernel.vhd:2557:104  */
  assign n5323_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:2557:95  */
  assign n5324_o = svmode | n5323_o;
  /* TG68KdotC_Kernel.vhd:2562:106  */
  assign n5326_o = opcode[2];
  assign n5329_o = n1909_o[59];
  /* TG68KdotC_Kernel.vhd:2562:97  */
  assign n5330_o = n5326_o ? n5329_o : 1'b1;
  assign n5331_o = n1909_o[60];
  /* TG68KdotC_Kernel.vhd:2562:97  */
  assign n5332_o = n5326_o ? 1'b1 : n5331_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5334_o = n5346_o ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5336_o = n5347_o ? 1'b1 : n2015_o;
  assign n5337_o = {n5332_o, n5330_o};
  assign n5338_o = n2162_o[0];
  assign n5339_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5340_o = n2037_o ? n5338_o : n5339_o;
  /* TG68KdotC_Kernel.vhd:2558:89  */
  assign n5341_o = decodeopc ? 1'b1 : n5340_o;
  assign n5342_o = n1909_o[60:59];
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5343_o = n5359_o ? n5337_o : n5342_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5345_o = n5360_o ? 7'b0101011 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5346_o = decodeopc & n5324_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5347_o = decodeopc & n5324_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5350_o = n5324_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5353_o = n5324_o ? 1'b0 : 1'b1;
  assign n5354_o = n2162_o[0];
  assign n5355_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5356_o = n2037_o ? n5354_o : n5355_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5357_o = n5324_o ? n5341_o : n5356_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5359_o = decodeopc & n5324_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5360_o = decodeopc & n5324_o;
  /* TG68KdotC_Kernel.vhd:2556:73  */
  assign n5362_o = n5061_o == 7'b1110011;
  /* TG68KdotC_Kernel.vhd:2556:87  */
  assign n5364_o = n5061_o == 7'b1110111;
  /* TG68KdotC_Kernel.vhd:2556:87  */
  assign n5365_o = n5362_o | n5364_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5370_o = decodeopc ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5372_o = decodeopc ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5374_o = decodeopc ? 1'b1 : n2154_o;
  assign n5375_o = {1'b1, 1'b1};
  assign n5376_o = n2162_o[0];
  assign n5377_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5378_o = n2037_o ? n5376_o : n5377_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5379_o = decodeopc ? 1'b1 : n5378_o;
  assign n5380_o = n1909_o[58:57];
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5381_o = decodeopc ? n5375_o : n5380_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5383_o = decodeopc ? 7'b0110000 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2574:73  */
  assign n5385_o = n5061_o == 7'b1110100;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5390_o = decodeopc ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5392_o = decodeopc ? 1'b1 : n2015_o;
  assign n5393_o = {1'b1, 1'b1};
  assign n5394_o = n2162_o[0];
  assign n5395_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5396_o = n2037_o ? n5394_o : n5395_o;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5397_o = decodeopc ? 1'b1 : n5396_o;
  assign n5398_o = n1909_o[58:57];
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5399_o = decodeopc ? n5393_o : n5398_o;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5401_o = decodeopc ? 7'b0011000 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2587:73  */
  assign n5403_o = n5061_o == 7'b1110101;
  /* TG68KdotC_Kernel.vhd:2599:81  */
  assign n5405_o = decodeopc ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2602:89  */
  assign n5406_o = flags[1];
  /* TG68KdotC_Kernel.vhd:2602:106  */
  assign n5408_o = state == 2'b01;
  /* TG68KdotC_Kernel.vhd:2602:97  */
  assign n5409_o = n5408_o & n5406_o;
  /* TG68KdotC_Kernel.vhd:2602:81  */
  assign n5412_o = n5409_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2602:81  */
  assign n5415_o = n5409_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2598:73  */
  assign n5417_o = n5061_o == 7'b1110110;
  /* TG68KdotC_Kernel.vhd:2608:87  */
  assign n5419_o = cpu == 2'b00;
  /* TG68KdotC_Kernel.vhd:2611:93  */
  assign n5420_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:2616:106  */
  assign n5421_o = last_data_read[11:0];
  /* TG68KdotC_Kernel.vhd:2616:119  */
  assign n5423_o = n5421_o == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:2618:106  */
  assign n5425_o = opcode[0];
  assign n5427_o = n2017_o[0];
  assign n5428_o = n1909_o[65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5429_o = n2010_o ? n5427_o : n5428_o;
  /* TG68KdotC_Kernel.vhd:2618:97  */
  assign n5430_o = n5425_o ? 1'b1 : n5429_o;
  assign n5431_o = {1'b1, n5430_o};
  /* TG68KdotC_Kernel.vhd:2616:89  */
  assign n5432_o = n5423_o ? n5431_o : n2019_o;
  /* TG68KdotC_Kernel.vhd:2622:98  */
  assign n5433_o = opcode[0];
  /* TG68KdotC_Kernel.vhd:2622:101  */
  assign n5434_o = ~n5433_o;
  /* TG68KdotC_Kernel.vhd:2622:89  */
  assign n5438_o = n5434_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2622:89  */
  assign n5440_o = n5434_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2627:89  */
  assign n5442_o = decodeopc ? 1'b1 : n2151_o;
  /* TG68KdotC_Kernel.vhd:2627:89  */
  assign n5444_o = decodeopc ? 7'b1001001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5446_o = n5420_o ? n1921_o : 2'b10;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5447_o = n5420_o ? n2151_o : n5442_o;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5450_o = n5420_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5453_o = n5420_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5454_o = n5420_o ? n2019_o : n5432_o;
  assign n5455_o = {n5440_o, n5438_o};
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5457_o = n5420_o ? 2'b00 : n5455_o;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5458_o = n5420_o ? n2180_o : n5444_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5459_o = n5419_o ? n1921_o : n5446_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5460_o = n5419_o ? n2151_o : n5447_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5463_o = n5419_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5465_o = n5419_o ? 1'b0 : n5450_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5467_o = n5419_o ? 1'b1 : n5453_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5468_o = n5419_o ? n2019_o : n5454_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5470_o = n5419_o ? 2'b00 : n5457_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5471_o = n5419_o ? n2180_o : n5458_o;
  /* TG68KdotC_Kernel.vhd:2607:73  */
  assign n5473_o = n5061_o == 7'b1111010;
  /* TG68KdotC_Kernel.vhd:2607:87  */
  assign n5475_o = n5061_o == 7'b1111011;
  /* TG68KdotC_Kernel.vhd:2607:87  */
  assign n5476_o = n5473_o | n5475_o;
  assign n5477_o = {n5476_o, n5417_o, n5403_o, n5385_o, n5365_o, n5322_o, n5302_o, n5300_o, n5280_o, n5241_o, n5199_o, n5155_o, n5108_o};
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5478_o = make_berr;
      13'b0100000000000: n5478_o = make_berr;
      13'b0010000000000: n5478_o = make_berr;
      13'b0001000000000: n5478_o = make_berr;
      13'b0000100000000: n5478_o = make_berr;
      13'b0000010000000: n5478_o = n5311_o;
      13'b0000001000000: n5478_o = make_berr;
      13'b0000000100000: n5478_o = make_berr;
      13'b0000000010000: n5478_o = make_berr;
      13'b0000000001000: n5478_o = make_berr;
      13'b0000000000100: n5478_o = make_berr;
      13'b0000000000010: n5478_o = make_berr;
      13'b0000000000001: n5478_o = make_berr;
      default: n5478_o = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5483_o = n5459_o;
      13'b0100000000000: n5483_o = n1921_o;
      13'b0010000000000: n5483_o = 2'b10;
      13'b0001000000000: n5483_o = 2'b10;
      13'b0000100000000: n5483_o = n1921_o;
      13'b0000010000000: n5483_o = n1921_o;
      13'b0000001000000: n5483_o = n1921_o;
      13'b0000000100000: n5483_o = n1921_o;
      13'b0000000010000: n5483_o = n5245_o;
      13'b0000000001000: n5483_o = n5202_o;
      13'b0000000000100: n5483_o = 2'b10;
      13'b0000000000010: n5483_o = 2'b10;
      13'b0000000000001: n5483_o = n1921_o;
      default: n5483_o = n1921_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5484_o = n2026_o;
      13'b0100000000000: n5484_o = n5405_o;
      13'b0010000000000: n5484_o = n5390_o;
      13'b0001000000000: n5484_o = n5370_o;
      13'b0000100000000: n5484_o = n5334_o;
      13'b0000010000000: n5484_o = n2026_o;
      13'b0000001000000: n5484_o = n2026_o;
      13'b0000000100000: n5484_o = n2026_o;
      13'b0000000010000: n5484_o = n2026_o;
      13'b0000000001000: n5484_o = n2026_o;
      13'b0000000000100: n5484_o = n5162_o;
      13'b0000000000010: n5484_o = n2026_o;
      13'b0000000000001: n5484_o = n2026_o;
      default: n5484_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5485_o = n2148_o;
      13'b0100000000000: n5485_o = n2148_o;
      13'b0010000000000: n5485_o = n2148_o;
      13'b0001000000000: n5485_o = n2148_o;
      13'b0000100000000: n5485_o = n2148_o;
      13'b0000010000000: n5485_o = n5312_o;
      13'b0000001000000: n5485_o = n2148_o;
      13'b0000000100000: n5485_o = n2148_o;
      13'b0000000010000: n5485_o = n2148_o;
      13'b0000000001000: n5485_o = n2148_o;
      13'b0000000000100: n5485_o = n2148_o;
      13'b0000000000010: n5485_o = n2148_o;
      13'b0000000000001: n5485_o = n2148_o;
      default: n5485_o = n2148_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5486_o = n5460_o;
      13'b0100000000000: n5486_o = n2151_o;
      13'b0010000000000: n5486_o = n2151_o;
      13'b0001000000000: n5486_o = n2151_o;
      13'b0000100000000: n5486_o = n2151_o;
      13'b0000010000000: n5486_o = n2151_o;
      13'b0000001000000: n5486_o = n2151_o;
      13'b0000000100000: n5486_o = n2151_o;
      13'b0000000010000: n5486_o = n2151_o;
      13'b0000000001000: n5486_o = n2151_o;
      13'b0000000000100: n5486_o = n2151_o;
      13'b0000000000010: n5486_o = n2151_o;
      13'b0000000000001: n5486_o = n2151_o;
      default: n5486_o = n2151_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5487_o = n2015_o;
      13'b0100000000000: n5487_o = n2015_o;
      13'b0010000000000: n5487_o = n5392_o;
      13'b0001000000000: n5487_o = n5372_o;
      13'b0000100000000: n5487_o = n5336_o;
      13'b0000010000000: n5487_o = n2015_o;
      13'b0000001000000: n5487_o = n2015_o;
      13'b0000000100000: n5487_o = n2015_o;
      13'b0000000010000: n5487_o = n2015_o;
      13'b0000000001000: n5487_o = n2015_o;
      13'b0000000000100: n5487_o = n5164_o;
      13'b0000000000010: n5487_o = n5116_o;
      13'b0000000000001: n5487_o = n2015_o;
      default: n5487_o = n2015_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5489_o = 1'b0;
      13'b0100000000000: n5489_o = 1'b0;
      13'b0010000000000: n5489_o = 1'b0;
      13'b0001000000000: n5489_o = 1'b0;
      13'b0000100000000: n5489_o = 1'b0;
      13'b0000010000000: n5489_o = 1'b0;
      13'b0000001000000: n5489_o = 1'b0;
      13'b0000000100000: n5489_o = 1'b0;
      13'b0000000010000: n5489_o = 1'b0;
      13'b0000000001000: n5489_o = n5205_o;
      13'b0000000000100: n5489_o = n5167_o;
      13'b0000000000010: n5489_o = n5119_o;
      13'b0000000000001: n5489_o = 1'b0;
      default: n5489_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5491_o = 1'b0;
      13'b0100000000000: n5491_o = 1'b0;
      13'b0010000000000: n5491_o = 1'b0;
      13'b0001000000000: n5491_o = 1'b0;
      13'b0000100000000: n5491_o = 1'b0;
      13'b0000010000000: n5491_o = 1'b0;
      13'b0000001000000: n5491_o = 1'b0;
      13'b0000000100000: n5491_o = 1'b0;
      13'b0000000010000: n5491_o = 1'b0;
      13'b0000000001000: n5491_o = n5208_o;
      13'b0000000000100: n5491_o = n5170_o;
      13'b0000000000010: n5491_o = n5122_o;
      13'b0000000000001: n5491_o = 1'b0;
      default: n5491_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5492_o = n1906_o;
      13'b0100000000000: n5492_o = n1906_o;
      13'b0010000000000: n5492_o = n1906_o;
      13'b0001000000000: n5492_o = n1906_o;
      13'b0000100000000: n5492_o = n1906_o;
      13'b0000010000000: n5492_o = n1906_o;
      13'b0000001000000: n5492_o = n1906_o;
      13'b0000000100000: n5492_o = n5288_o;
      13'b0000000010000: n5492_o = n1906_o;
      13'b0000000001000: n5492_o = n1906_o;
      13'b0000000000100: n5492_o = n1906_o;
      13'b0000000000010: n5492_o = n1906_o;
      13'b0000000000001: n5492_o = n1906_o;
      default: n5492_o = n1906_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5493_o = n2154_o;
      13'b0100000000000: n5493_o = n2154_o;
      13'b0010000000000: n5493_o = n2154_o;
      13'b0001000000000: n5493_o = n5374_o;
      13'b0000100000000: n5493_o = n2154_o;
      13'b0000010000000: n5493_o = n2154_o;
      13'b0000001000000: n5493_o = n2154_o;
      13'b0000000100000: n5493_o = n2154_o;
      13'b0000000010000: n5493_o = n2154_o;
      13'b0000000001000: n5493_o = n2154_o;
      13'b0000000000100: n5493_o = n2154_o;
      13'b0000000000010: n5493_o = n2154_o;
      13'b0000000000001: n5493_o = n2154_o;
      default: n5493_o = n2154_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5496_o = n5463_o;
      13'b0100000000000: n5496_o = 1'b0;
      13'b0010000000000: n5496_o = 1'b0;
      13'b0001000000000: n5496_o = 1'b0;
      13'b0000100000000: n5496_o = 1'b0;
      13'b0000010000000: n5496_o = 1'b0;
      13'b0000001000000: n5496_o = 1'b0;
      13'b0000000100000: n5496_o = 1'b0;
      13'b0000000010000: n5496_o = 1'b0;
      13'b0000000001000: n5496_o = 1'b0;
      13'b0000000000100: n5496_o = 1'b0;
      13'b0000000000010: n5496_o = 1'b0;
      13'b0000000000001: n5496_o = 1'b0;
      default: n5496_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5498_o = n5465_o;
      13'b0100000000000: n5498_o = 1'b0;
      13'b0010000000000: n5498_o = 1'b0;
      13'b0001000000000: n5498_o = 1'b0;
      13'b0000100000000: n5498_o = n5350_o;
      13'b0000010000000: n5498_o = n5315_o;
      13'b0000001000000: n5498_o = 1'b0;
      13'b0000000100000: n5498_o = n5291_o;
      13'b0000000010000: n5498_o = n5248_o;
      13'b0000000001000: n5498_o = n5211_o;
      13'b0000000000100: n5498_o = 1'b0;
      13'b0000000000010: n5498_o = 1'b0;
      13'b0000000000001: n5498_o = 1'b0;
      default: n5498_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5501_o = 1'b0;
      13'b0100000000000: n5501_o = 1'b0;
      13'b0010000000000: n5501_o = 1'b0;
      13'b0001000000000: n5501_o = 1'b0;
      13'b0000100000000: n5501_o = 1'b0;
      13'b0000010000000: n5501_o = 1'b0;
      13'b0000001000000: n5501_o = 1'b0;
      13'b0000000100000: n5501_o = 1'b0;
      13'b0000000010000: n5501_o = 1'b0;
      13'b0000000001000: n5501_o = 1'b0;
      13'b0000000000100: n5501_o = 1'b0;
      13'b0000000000010: n5501_o = 1'b0;
      13'b0000000000001: n5501_o = 1'b1;
      default: n5501_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5503_o = 1'b0;
      13'b0100000000000: n5503_o = n5412_o;
      13'b0010000000000: n5503_o = 1'b0;
      13'b0001000000000: n5503_o = 1'b0;
      13'b0000100000000: n5503_o = 1'b0;
      13'b0000010000000: n5503_o = 1'b0;
      13'b0000001000000: n5503_o = 1'b0;
      13'b0000000100000: n5503_o = 1'b0;
      13'b0000000010000: n5503_o = 1'b0;
      13'b0000000001000: n5503_o = 1'b0;
      13'b0000000000100: n5503_o = 1'b0;
      13'b0000000000010: n5503_o = 1'b0;
      13'b0000000000001: n5503_o = 1'b0;
      default: n5503_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5507_o = n5467_o;
      13'b0100000000000: n5507_o = n5415_o;
      13'b0010000000000: n5507_o = 1'b0;
      13'b0001000000000: n5507_o = 1'b0;
      13'b0000100000000: n5507_o = n5353_o;
      13'b0000010000000: n5507_o = n5318_o;
      13'b0000001000000: n5507_o = 1'b0;
      13'b0000000100000: n5507_o = n5294_o;
      13'b0000000010000: n5507_o = n5251_o;
      13'b0000000001000: n5507_o = n5214_o;
      13'b0000000000100: n5507_o = 1'b0;
      13'b0000000000010: n5507_o = 1'b0;
      13'b0000000000001: n5507_o = 1'b1;
      default: n5507_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5509_o = 1'b0;
      13'b0100000000000: n5509_o = 1'b0;
      13'b0010000000000: n5509_o = 1'b0;
      13'b0001000000000: n5509_o = 1'b0;
      13'b0000100000000: n5509_o = 1'b0;
      13'b0000010000000: n5509_o = n5320_o;
      13'b0000001000000: n5509_o = 1'b0;
      13'b0000000100000: n5509_o = 1'b0;
      13'b0000000010000: n5509_o = 1'b0;
      13'b0000000001000: n5509_o = 1'b0;
      13'b0000000000100: n5509_o = 1'b0;
      13'b0000000000010: n5509_o = 1'b0;
      13'b0000000000001: n5509_o = 1'b0;
      default: n5509_o = 1'b0;
    endcase
  assign n5510_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5511_o = n5510_o;
      13'b0100000000000: n5511_o = n5510_o;
      13'b0010000000000: n5511_o = n5510_o;
      13'b0001000000000: n5511_o = n5510_o;
      13'b0000100000000: n5511_o = n5510_o;
      13'b0000010000000: n5511_o = n5510_o;
      13'b0000001000000: n5511_o = n5510_o;
      13'b0000000100000: n5511_o = n5510_o;
      13'b0000000010000: n5511_o = n5510_o;
      13'b0000000001000: n5511_o = n5510_o;
      13'b0000000000100: n5511_o = n5172_o;
      13'b0000000000010: n5511_o = n5510_o;
      13'b0000000000001: n5511_o = n5510_o;
      default: n5511_o = n5510_o;
    endcase
  assign n5512_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5513_o = n5512_o;
      13'b0100000000000: n5513_o = n5512_o;
      13'b0010000000000: n5513_o = n5512_o;
      13'b0001000000000: n5513_o = n5512_o;
      13'b0000100000000: n5513_o = n5512_o;
      13'b0000010000000: n5513_o = n5512_o;
      13'b0000001000000: n5513_o = n5512_o;
      13'b0000000100000: n5513_o = n5296_o;
      13'b0000000010000: n5513_o = n5512_o;
      13'b0000000001000: n5513_o = n5512_o;
      13'b0000000000100: n5513_o = n5512_o;
      13'b0000000000010: n5513_o = n5512_o;
      13'b0000000000001: n5513_o = n5512_o;
      default: n5513_o = n5512_o;
    endcase
  assign n5514_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5515_o = n5514_o;
      13'b0100000000000: n5515_o = n5514_o;
      13'b0010000000000: n5515_o = n5514_o;
      13'b0001000000000: n5515_o = n5514_o;
      13'b0000100000000: n5515_o = n5514_o;
      13'b0000010000000: n5515_o = n5514_o;
      13'b0000001000000: n5515_o = n5514_o;
      13'b0000000100000: n5515_o = n5514_o;
      13'b0000000010000: n5515_o = n5514_o;
      13'b0000000001000: n5515_o = n5514_o;
      13'b0000000000100: n5515_o = n5174_o;
      13'b0000000000010: n5515_o = n5514_o;
      13'b0000000000001: n5515_o = n5514_o;
      default: n5515_o = n5514_o;
    endcase
  assign n5516_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5517_o = n5516_o;
      13'b0100000000000: n5517_o = n5516_o;
      13'b0010000000000: n5517_o = n5516_o;
      13'b0001000000000: n5517_o = n5516_o;
      13'b0000100000000: n5517_o = n5516_o;
      13'b0000010000000: n5517_o = n5516_o;
      13'b0000001000000: n5517_o = n5516_o;
      13'b0000000100000: n5517_o = n5516_o;
      13'b0000000010000: n5517_o = n5516_o;
      13'b0000000001000: n5517_o = n5516_o;
      13'b0000000000100: n5517_o = n5516_o;
      13'b0000000000010: n5517_o = n5124_o;
      13'b0000000000001: n5517_o = n5516_o;
      default: n5517_o = n5516_o;
    endcase
  assign n5518_o = n2162_o[0];
  assign n5519_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5520_o = n2037_o ? n5518_o : n5519_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5521_o = n5520_o;
      13'b0100000000000: n5521_o = n5520_o;
      13'b0010000000000: n5521_o = n5397_o;
      13'b0001000000000: n5521_o = n5379_o;
      13'b0000100000000: n5521_o = n5357_o;
      13'b0000010000000: n5521_o = n5520_o;
      13'b0000001000000: n5521_o = n5520_o;
      13'b0000000100000: n5521_o = n5520_o;
      13'b0000000010000: n5521_o = n5520_o;
      13'b0000000001000: n5521_o = n5520_o;
      13'b0000000000100: n5521_o = n5520_o;
      13'b0000000000010: n5521_o = n5520_o;
      13'b0000000000001: n5521_o = n5520_o;
      default: n5521_o = n5520_o;
    endcase
  assign n5522_o = n2162_o[1];
  assign n5523_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5524_o = n2037_o ? n5522_o : n5523_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5525_o = n5524_o;
      13'b0100000000000: n5525_o = n5524_o;
      13'b0010000000000: n5525_o = n5524_o;
      13'b0001000000000: n5525_o = n5524_o;
      13'b0000100000000: n5525_o = n5524_o;
      13'b0000010000000: n5525_o = n5524_o;
      13'b0000001000000: n5525_o = n5524_o;
      13'b0000000100000: n5525_o = n5524_o;
      13'b0000000010000: n5525_o = n5524_o;
      13'b0000000001000: n5525_o = n5524_o;
      13'b0000000000100: n5525_o = n5524_o;
      13'b0000000000010: n5525_o = n5128_o;
      13'b0000000000001: n5525_o = n5524_o;
      default: n5525_o = n5524_o;
    endcase
  assign n5526_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5527_o = n5526_o;
      13'b0100000000000: n5527_o = n5526_o;
      13'b0010000000000: n5527_o = n5526_o;
      13'b0001000000000: n5527_o = n5526_o;
      13'b0000100000000: n5527_o = n5526_o;
      13'b0000010000000: n5527_o = n5526_o;
      13'b0000001000000: n5527_o = n5526_o;
      13'b0000000100000: n5527_o = n5526_o;
      13'b0000000010000: n5527_o = n5526_o;
      13'b0000000001000: n5527_o = n5526_o;
      13'b0000000000100: n5527_o = 1'b1;
      13'b0000000000010: n5527_o = 1'b1;
      13'b0000000000001: n5527_o = n5526_o;
      default: n5527_o = n5526_o;
    endcase
  assign n5528_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5529_o = n5528_o;
      13'b0100000000000: n5529_o = n5528_o;
      13'b0010000000000: n5529_o = n5528_o;
      13'b0001000000000: n5529_o = n5528_o;
      13'b0000100000000: n5529_o = n5528_o;
      13'b0000010000000: n5529_o = n5528_o;
      13'b0000001000000: n5529_o = n5528_o;
      13'b0000000100000: n5529_o = n5528_o;
      13'b0000000010000: n5529_o = n5528_o;
      13'b0000000001000: n5529_o = n5528_o;
      13'b0000000000100: n5529_o = n5528_o;
      13'b0000000000010: n5529_o = n5130_o;
      13'b0000000000001: n5529_o = n5528_o;
      default: n5529_o = n5528_o;
    endcase
  assign n5530_o = n1909_o[58:57];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5531_o = n5530_o;
      13'b0100000000000: n5531_o = n5530_o;
      13'b0010000000000: n5531_o = n5399_o;
      13'b0001000000000: n5531_o = n5381_o;
      13'b0000100000000: n5531_o = n5530_o;
      13'b0000010000000: n5531_o = n5530_o;
      13'b0000001000000: n5531_o = n5530_o;
      13'b0000000100000: n5531_o = n5530_o;
      13'b0000000010000: n5531_o = n5530_o;
      13'b0000000001000: n5531_o = n5530_o;
      13'b0000000000100: n5531_o = n5530_o;
      13'b0000000000010: n5531_o = n5530_o;
      13'b0000000000001: n5531_o = n5530_o;
      default: n5531_o = n5530_o;
    endcase
  assign n5532_o = n1909_o[60:59];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5533_o = n5532_o;
      13'b0100000000000: n5533_o = n5532_o;
      13'b0010000000000: n5533_o = n5532_o;
      13'b0001000000000: n5533_o = n5532_o;
      13'b0000100000000: n5533_o = n5343_o;
      13'b0000010000000: n5533_o = n5532_o;
      13'b0000001000000: n5533_o = n5532_o;
      13'b0000000100000: n5533_o = n5532_o;
      13'b0000000010000: n5533_o = n5532_o;
      13'b0000000001000: n5533_o = n5532_o;
      13'b0000000000100: n5533_o = n5532_o;
      13'b0000000000010: n5533_o = n5532_o;
      13'b0000000000001: n5533_o = n5532_o;
      default: n5533_o = n5532_o;
    endcase
  assign n5534_o = n5468_o[0];
  assign n5535_o = n2017_o[0];
  assign n5536_o = n1909_o[65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5537_o = n2010_o ? n5535_o : n5536_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5538_o = n5534_o;
      13'b0100000000000: n5538_o = n5537_o;
      13'b0010000000000: n5538_o = n5537_o;
      13'b0001000000000: n5538_o = n5537_o;
      13'b0000100000000: n5538_o = n5537_o;
      13'b0000010000000: n5538_o = n5537_o;
      13'b0000001000000: n5538_o = n5537_o;
      13'b0000000100000: n5538_o = n5537_o;
      13'b0000000010000: n5538_o = n5537_o;
      13'b0000000001000: n5538_o = n5218_o;
      13'b0000000000100: n5538_o = n5537_o;
      13'b0000000000010: n5538_o = n5537_o;
      13'b0000000000001: n5538_o = n5537_o;
      default: n5538_o = n5537_o;
    endcase
  assign n5539_o = n5468_o[1];
  assign n5540_o = n2017_o[1];
  assign n5541_o = n1909_o[66];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5542_o = n2010_o ? n5540_o : n5541_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5543_o = n5539_o;
      13'b0100000000000: n5543_o = n5542_o;
      13'b0010000000000: n5543_o = n5542_o;
      13'b0001000000000: n5543_o = n5542_o;
      13'b0000100000000: n5543_o = n5542_o;
      13'b0000010000000: n5543_o = n5542_o;
      13'b0000001000000: n5543_o = n5542_o;
      13'b0000000100000: n5543_o = n5542_o;
      13'b0000000010000: n5543_o = n5255_o;
      13'b0000000001000: n5543_o = n5542_o;
      13'b0000000000100: n5543_o = n5542_o;
      13'b0000000000010: n5543_o = n5542_o;
      13'b0000000000001: n5543_o = n5542_o;
      default: n5543_o = n5542_o;
    endcase
  assign n5544_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5545_o = n5544_o;
      13'b0100000000000: n5545_o = n5544_o;
      13'b0010000000000: n5545_o = n5544_o;
      13'b0001000000000: n5545_o = n5544_o;
      13'b0000100000000: n5545_o = n5544_o;
      13'b0000010000000: n5545_o = n5544_o;
      13'b0000001000000: n5545_o = n5544_o;
      13'b0000000100000: n5545_o = n5298_o;
      13'b0000000010000: n5545_o = n5544_o;
      13'b0000000001000: n5545_o = n5544_o;
      13'b0000000000100: n5545_o = n5544_o;
      13'b0000000000010: n5545_o = n5544_o;
      13'b0000000000001: n5545_o = n5544_o;
      default: n5545_o = n5544_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5547_o = 1'b0;
      13'b0100000000000: n5547_o = 1'b0;
      13'b0010000000000: n5547_o = 1'b0;
      13'b0001000000000: n5547_o = 1'b0;
      13'b0000100000000: n5547_o = 1'b0;
      13'b0000010000000: n5547_o = 1'b0;
      13'b0000001000000: n5547_o = 1'b0;
      13'b0000000100000: n5547_o = 1'b0;
      13'b0000000010000: n5547_o = 1'b0;
      13'b0000000001000: n5547_o = 1'b0;
      13'b0000000000100: n5547_o = 1'b1;
      13'b0000000000010: n5547_o = 1'b0;
      13'b0000000000001: n5547_o = 1'b0;
      default: n5547_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5549_o = 1'b0;
      13'b0100000000000: n5549_o = 1'b0;
      13'b0010000000000: n5549_o = 1'b0;
      13'b0001000000000: n5549_o = 1'b0;
      13'b0000100000000: n5549_o = 1'b0;
      13'b0000010000000: n5549_o = 1'b0;
      13'b0000001000000: n5549_o = 1'b0;
      13'b0000000100000: n5549_o = 1'b0;
      13'b0000000010000: n5549_o = 1'b0;
      13'b0000000001000: n5549_o = 1'b0;
      13'b0000000000100: n5549_o = 1'b0;
      13'b0000000000010: n5549_o = 1'b1;
      13'b0000000000001: n5549_o = 1'b0;
      default: n5549_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5551_o = n5470_o;
      13'b0100000000000: n5551_o = 2'b00;
      13'b0010000000000: n5551_o = 2'b00;
      13'b0001000000000: n5551_o = 2'b00;
      13'b0000100000000: n5551_o = 2'b00;
      13'b0000010000000: n5551_o = 2'b00;
      13'b0000001000000: n5551_o = 2'b00;
      13'b0000000100000: n5551_o = 2'b00;
      13'b0000000010000: n5551_o = 2'b00;
      13'b0000000001000: n5551_o = 2'b00;
      13'b0000000000100: n5551_o = 2'b00;
      13'b0000000000010: n5551_o = 2'b00;
      13'b0000000000001: n5551_o = 2'b00;
      default: n5551_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5553_o = 1'b0;
      13'b0100000000000: n5553_o = 1'b0;
      13'b0010000000000: n5553_o = 1'b0;
      13'b0001000000000: n5553_o = 1'b0;
      13'b0000100000000: n5553_o = 1'b0;
      13'b0000010000000: n5553_o = 1'b0;
      13'b0000001000000: n5553_o = 1'b0;
      13'b0000000100000: n5553_o = 1'b0;
      13'b0000000010000: n5553_o = n5257_o;
      13'b0000000001000: n5553_o = 1'b0;
      13'b0000000000100: n5553_o = 1'b1;
      13'b0000000000010: n5553_o = 1'b1;
      13'b0000000000001: n5553_o = 1'b0;
      default: n5553_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5477_o)
      13'b1000000000000: n5554_o = n5471_o;
      13'b0100000000000: n5554_o = n2180_o;
      13'b0010000000000: n5554_o = n5401_o;
      13'b0001000000000: n5554_o = n5383_o;
      13'b0000100000000: n5554_o = n5345_o;
      13'b0000010000000: n5554_o = n2180_o;
      13'b0000001000000: n5554_o = n2180_o;
      13'b0000000100000: n5554_o = n2180_o;
      13'b0000000010000: n5554_o = n2180_o;
      13'b0000000001000: n5554_o = n2180_o;
      13'b0000000000100: n5554_o = n5176_o;
      13'b0000000000010: n5554_o = n5132_o;
      13'b0000000000001: n5554_o = n2180_o;
      default: n5554_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5555_o = n4976_o ? n5035_o : n5478_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5556_o = n4976_o ? n5037_o : n5483_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5557_o = n4976_o ? n5038_o : n5484_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5558_o = n4976_o ? n2148_o : n5485_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5559_o = n4976_o ? n2151_o : n5486_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5560_o = n4976_o ? n5003_o : n5487_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5562_o = n4976_o ? n5041_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5564_o = n4976_o ? n5044_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5566_o = n4976_o ? 1'b0 : n5489_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5568_o = n4976_o ? 1'b0 : n5491_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5569_o = n4976_o ? n1906_o : n5492_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5570_o = n4976_o ? n2154_o : n5493_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5571_o = n4976_o ? n5047_o : n5496_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5573_o = n4976_o ? 1'b0 : n5498_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5575_o = n4976_o ? 1'b0 : n5501_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5577_o = n4976_o ? 1'b0 : n5503_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5578_o = n4976_o ? n5050_o : n5507_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5580_o = n4976_o ? 1'b0 : n5509_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5582_o = n4976_o ? n5053_o : 1'b0;
  assign n5583_o = {n5525_o, n5521_o};
  assign n5584_o = {n5533_o, n5531_o};
  assign n5585_o = {n5543_o, n5538_o};
  assign n5586_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5587_o = n4976_o ? n5586_o : n5511_o;
  assign n5588_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5589_o = n4976_o ? n5588_o : n5513_o;
  assign n5590_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5591_o = n4976_o ? n5590_o : n5515_o;
  assign n5592_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5593_o = n4976_o ? n5592_o : n5517_o;
  assign n5594_o = n5583_o[0];
  assign n5595_o = n2162_o[0];
  assign n5596_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5597_o = n2037_o ? n5595_o : n5596_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5598_o = n4976_o ? n5597_o : n5594_o;
  assign n5599_o = n5583_o[1];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5600_o = n4976_o ? n5058_o : n5599_o;
  assign n5601_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5602_o = n4976_o ? n5601_o : n5527_o;
  assign n5603_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5604_o = n4976_o ? n5603_o : n5529_o;
  assign n5605_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5606_o = n4976_o ? n5605_o : n5584_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5607_o = n4989_o & n4976_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5608_o = n4976_o ? n2019_o : n5585_o;
  assign n5609_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5610_o = n4976_o ? n5609_o : n5545_o;
  assign n5611_o = {n5553_o, n5551_o};
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5613_o = n4976_o ? 1'b0 : n5547_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5615_o = n4976_o ? 1'b0 : n5549_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5617_o = n4976_o ? 3'b000 : n5611_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5618_o = n4976_o ? n5060_o : n5554_o;
  /* TG68KdotC_Kernel.vhd:2415:49  */
  assign n5620_o = n3613_o == 3'b111;
  assign n5621_o = {n5620_o, n4975_o, n4865_o, n4078_o, n3938_o, n3831_o, n3732_o};
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5622_o = n5555_o;
      7'b0100000: n5622_o = make_berr;
      7'b0010000: n5622_o = make_berr;
      7'b0001000: n5622_o = make_berr;
      7'b0000100: n5622_o = make_berr;
      7'b0000010: n5622_o = n3812_o;
      7'b0000001: n5622_o = n3643_o;
      default: n5622_o = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5623_o = n5556_o;
      7'b0100000: n5623_o = n4955_o;
      7'b0010000: n5623_o = n4785_o;
      7'b0001000: n5623_o = n3983_o;
      7'b0000100: n5623_o = n3860_o;
      7'b0000010: n5623_o = n3760_o;
      7'b0000001: n5623_o = n3652_o;
      default: n5623_o = n1921_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5624_o = n5557_o;
      7'b0100000: n5624_o = n2026_o;
      7'b0010000: n5624_o = n4786_o;
      7'b0001000: n5624_o = n3981_o;
      7'b0000100: n5624_o = n2026_o;
      7'b0000010: n5624_o = n2026_o;
      7'b0000001: n5624_o = n2026_o;
      default: n5624_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5625_o = n5558_o;
      7'b0100000: n5625_o = n2148_o;
      7'b0010000: n5625_o = n2148_o;
      7'b0001000: n5625_o = n2148_o;
      7'b0000100: n5625_o = n2148_o;
      7'b0000010: n5625_o = n2148_o;
      7'b0000001: n5625_o = n2148_o;
      default: n5625_o = n2148_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5626_o = n5559_o;
      7'b0100000: n5626_o = n2151_o;
      7'b0010000: n5626_o = n2151_o;
      7'b0001000: n5626_o = n2151_o;
      7'b0000100: n5626_o = n2151_o;
      7'b0000010: n5626_o = n2151_o;
      7'b0000001: n5626_o = n2151_o;
      default: n5626_o = n2151_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5628_o = 1'b0;
      7'b0100000: n5628_o = n4957_o;
      7'b0010000: n5628_o = n4788_o;
      7'b0001000: n5628_o = n4059_o;
      7'b0000100: n5628_o = n3922_o;
      7'b0000010: n5628_o = n3815_o;
      7'b0000001: n5628_o = n3708_o;
      default: n5628_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5629_o = n5560_o;
      7'b0100000: n5629_o = n2015_o;
      7'b0010000: n5629_o = n4789_o;
      7'b0001000: n5629_o = n2015_o;
      7'b0000100: n5629_o = n2015_o;
      7'b0000010: n5629_o = n2015_o;
      7'b0000001: n5629_o = n2015_o;
      default: n5629_o = n2015_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5631_o = n5562_o;
      7'b0100000: n5631_o = 1'b0;
      7'b0010000: n5631_o = 1'b0;
      7'b0001000: n5631_o = 1'b0;
      7'b0000100: n5631_o = 1'b0;
      7'b0000010: n5631_o = 1'b0;
      7'b0000001: n5631_o = 1'b0;
      default: n5631_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5633_o = 1'b0;
      7'b0100000: n5633_o = n4959_o;
      7'b0010000: n5633_o = 1'b0;
      7'b0001000: n5633_o = 1'b0;
      7'b0000100: n5633_o = 1'b0;
      7'b0000010: n5633_o = 1'b0;
      7'b0000001: n5633_o = 1'b0;
      default: n5633_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5635_o = n5564_o;
      7'b0100000: n5635_o = 1'b0;
      7'b0010000: n5635_o = n4790_o;
      7'b0001000: n5635_o = 1'b0;
      7'b0000100: n5635_o = 1'b0;
      7'b0000010: n5635_o = 1'b0;
      7'b0000001: n5635_o = 1'b0;
      default: n5635_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5637_o = n5566_o;
      7'b0100000: n5637_o = n4961_o;
      7'b0010000: n5637_o = n4792_o;
      7'b0001000: n5637_o = 1'b0;
      7'b0000100: n5637_o = 1'b0;
      7'b0000010: n5637_o = 1'b0;
      7'b0000001: n5637_o = 1'b0;
      default: n5637_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5639_o = n5568_o;
      7'b0100000: n5639_o = n4963_o;
      7'b0010000: n5639_o = n4793_o;
      7'b0001000: n5639_o = n4061_o;
      7'b0000100: n5639_o = n3923_o;
      7'b0000010: n5639_o = 1'b0;
      7'b0000001: n5639_o = n3710_o;
      default: n5639_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5641_o = 1'b0;
      7'b0100000: n5641_o = 1'b0;
      7'b0010000: n5641_o = n4795_o;
      7'b0001000: n5641_o = 1'b0;
      7'b0000100: n5641_o = 1'b0;
      7'b0000010: n5641_o = 1'b0;
      7'b0000001: n5641_o = 1'b0;
      default: n5641_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5643_o = 1'b0;
      7'b0100000: n5643_o = 1'b0;
      7'b0010000: n5643_o = n4797_o;
      7'b0001000: n5643_o = 1'b0;
      7'b0000100: n5643_o = 1'b0;
      7'b0000010: n5643_o = 1'b0;
      7'b0000001: n5643_o = 1'b0;
      default: n5643_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5645_o = 1'b0;
      7'b0100000: n5645_o = 1'b0;
      7'b0010000: n5645_o = n4799_o;
      7'b0001000: n5645_o = 1'b0;
      7'b0000100: n5645_o = 1'b0;
      7'b0000010: n5645_o = 1'b0;
      7'b0000001: n5645_o = 1'b0;
      default: n5645_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5646_o = n5569_o;
      7'b0100000: n5646_o = n1906_o;
      7'b0010000: n5646_o = n1906_o;
      7'b0001000: n5646_o = n1906_o;
      7'b0000100: n5646_o = n1906_o;
      7'b0000010: n5646_o = n1906_o;
      7'b0000001: n5646_o = n1906_o;
      default: n5646_o = n1906_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5648_o = 1'b0;
      7'b0100000: n5648_o = 1'b0;
      7'b0010000: n5648_o = n4801_o;
      7'b0001000: n5648_o = 1'b0;
      7'b0000100: n5648_o = 1'b0;
      7'b0000010: n5648_o = 1'b0;
      7'b0000001: n5648_o = 1'b0;
      default: n5648_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5649_o = n5570_o;
      7'b0100000: n5649_o = n2154_o;
      7'b0010000: n5649_o = n2154_o;
      7'b0001000: n5649_o = n2154_o;
      7'b0000100: n5649_o = n2154_o;
      7'b0000010: n5649_o = n2154_o;
      7'b0000001: n5649_o = n2154_o;
      default: n5649_o = n2154_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5651_o = n5571_o;
      7'b0100000: n5651_o = n4965_o;
      7'b0010000: n5651_o = n4802_o;
      7'b0001000: n5651_o = n4062_o;
      7'b0000100: n5651_o = n3924_o;
      7'b0000010: n5651_o = n3817_o;
      7'b0000001: n5651_o = n3713_o;
      default: n5651_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5653_o = n5573_o;
      7'b0100000: n5653_o = 1'b0;
      7'b0010000: n5653_o = 1'b0;
      7'b0001000: n5653_o = n4064_o;
      7'b0000100: n5653_o = 1'b0;
      7'b0000010: n5653_o = 1'b0;
      7'b0000001: n5653_o = n3715_o;
      default: n5653_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5655_o = n5575_o;
      7'b0100000: n5655_o = 1'b0;
      7'b0010000: n5655_o = 1'b0;
      7'b0001000: n5655_o = 1'b0;
      7'b0000100: n5655_o = 1'b0;
      7'b0000010: n5655_o = 1'b0;
      7'b0000001: n5655_o = 1'b0;
      default: n5655_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5657_o = n5577_o;
      7'b0100000: n5657_o = 1'b0;
      7'b0010000: n5657_o = 1'b0;
      7'b0001000: n5657_o = 1'b0;
      7'b0000100: n5657_o = 1'b0;
      7'b0000010: n5657_o = 1'b0;
      7'b0000001: n5657_o = 1'b0;
      default: n5657_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5659_o = n5578_o;
      7'b0100000: n5659_o = n4967_o;
      7'b0010000: n5659_o = n4803_o;
      7'b0001000: n5659_o = n4065_o;
      7'b0000100: n5659_o = n3925_o;
      7'b0000010: n5659_o = n3819_o;
      7'b0000001: n5659_o = n3717_o;
      default: n5659_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5661_o = n5580_o;
      7'b0100000: n5661_o = 1'b0;
      7'b0010000: n5661_o = 1'b0;
      7'b0001000: n5661_o = 1'b0;
      7'b0000100: n5661_o = 1'b0;
      7'b0000010: n5661_o = 1'b0;
      7'b0000001: n5661_o = 1'b0;
      default: n5661_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5663_o = n5582_o;
      7'b0100000: n5663_o = n4969_o;
      7'b0010000: n5663_o = n4805_o;
      7'b0001000: n5663_o = n4066_o;
      7'b0000100: n5663_o = n3926_o;
      7'b0000010: n5663_o = n3821_o;
      7'b0000001: n5663_o = n3719_o;
      default: n5663_o = 1'b0;
    endcase
  assign n5664_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5665_o = n5587_o;
      7'b0100000: n5665_o = n5664_o;
      7'b0010000: n5665_o = n4807_o;
      7'b0001000: n5665_o = n5664_o;
      7'b0000100: n5665_o = n5664_o;
      7'b0000010: n5665_o = n5664_o;
      7'b0000001: n5665_o = n5664_o;
      default: n5665_o = n5664_o;
    endcase
  assign n5666_o = n1909_o[20];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5667_o = n5666_o;
      7'b0100000: n5667_o = n5666_o;
      7'b0010000: n5667_o = n4809_o;
      7'b0001000: n5667_o = n5666_o;
      7'b0000100: n5667_o = n5666_o;
      7'b0000010: n5667_o = n5666_o;
      7'b0000001: n5667_o = n5666_o;
      default: n5667_o = n5666_o;
    endcase
  assign n5668_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5669_o = n5589_o;
      7'b0100000: n5669_o = n5668_o;
      7'b0010000: n5669_o = n4811_o;
      7'b0001000: n5669_o = n5668_o;
      7'b0000100: n5669_o = n5668_o;
      7'b0000010: n5669_o = n5668_o;
      7'b0000001: n5669_o = n5668_o;
      default: n5669_o = n5668_o;
    endcase
  assign n5670_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5671_o = n5591_o;
      7'b0100000: n5671_o = n5670_o;
      7'b0010000: n5671_o = n4812_o;
      7'b0001000: n5671_o = n5670_o;
      7'b0000100: n5671_o = n5670_o;
      7'b0000010: n5671_o = n5670_o;
      7'b0000001: n5671_o = n5670_o;
      default: n5671_o = n5670_o;
    endcase
  assign n5672_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5673_o = n5672_o;
      7'b0100000: n5673_o = n5672_o;
      7'b0010000: n5673_o = n4814_o;
      7'b0001000: n5673_o = n5672_o;
      7'b0000100: n5673_o = n5672_o;
      7'b0000010: n5673_o = n5672_o;
      7'b0000001: n5673_o = n5672_o;
      default: n5673_o = n5672_o;
    endcase
  assign n5674_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5675_o = n5674_o;
      7'b0100000: n5675_o = n5674_o;
      7'b0010000: n5675_o = n4816_o;
      7'b0001000: n5675_o = n5674_o;
      7'b0000100: n5675_o = n5674_o;
      7'b0000010: n5675_o = n5674_o;
      7'b0000001: n5675_o = n5674_o;
      default: n5675_o = n5674_o;
    endcase
  assign n5676_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5677_o = n5676_o;
      7'b0100000: n5677_o = n5676_o;
      7'b0010000: n5677_o = n4817_o;
      7'b0001000: n5677_o = n5676_o;
      7'b0000100: n5677_o = n5676_o;
      7'b0000010: n5677_o = n5676_o;
      7'b0000001: n5677_o = n5676_o;
      default: n5677_o = n5676_o;
    endcase
  assign n5678_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5679_o = n5593_o;
      7'b0100000: n5679_o = n5678_o;
      7'b0010000: n5679_o = n4819_o;
      7'b0001000: n5679_o = n5678_o;
      7'b0000100: n5679_o = n5678_o;
      7'b0000010: n5679_o = n5678_o;
      7'b0000001: n5679_o = n5678_o;
      default: n5679_o = n5678_o;
    endcase
  assign n5680_o = n2162_o[0];
  assign n5681_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5682_o = n2037_o ? n5680_o : n5681_o;
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5683_o = n5598_o;
      7'b0100000: n5683_o = n5682_o;
      7'b0010000: n5683_o = n5682_o;
      7'b0001000: n5683_o = n5682_o;
      7'b0000100: n5683_o = n5682_o;
      7'b0000010: n5683_o = n5682_o;
      7'b0000001: n5683_o = n5682_o;
      default: n5683_o = n5682_o;
    endcase
  assign n5684_o = n2162_o[1];
  assign n5685_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5686_o = n2037_o ? n5684_o : n5685_o;
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5687_o = n5600_o;
      7'b0100000: n5687_o = n5686_o;
      7'b0010000: n5687_o = n4823_o;
      7'b0001000: n5687_o = n5686_o;
      7'b0000100: n5687_o = n5686_o;
      7'b0000010: n5687_o = n5686_o;
      7'b0000001: n5687_o = n5686_o;
      default: n5687_o = n5686_o;
    endcase
  assign n5688_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5689_o = n5688_o;
      7'b0100000: n5689_o = n5688_o;
      7'b0010000: n5689_o = n4826_o;
      7'b0001000: n5689_o = n5688_o;
      7'b0000100: n5689_o = n5688_o;
      7'b0000010: n5689_o = n5688_o;
      7'b0000001: n5689_o = n5688_o;
      default: n5689_o = n5688_o;
    endcase
  assign n5690_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5691_o = n5602_o;
      7'b0100000: n5691_o = n5690_o;
      7'b0010000: n5691_o = n4828_o;
      7'b0001000: n5691_o = n5690_o;
      7'b0000100: n5691_o = n5690_o;
      7'b0000010: n5691_o = n5690_o;
      7'b0000001: n5691_o = n5690_o;
      default: n5691_o = n5690_o;
    endcase
  assign n5692_o = n3967_o[0];
  assign n5693_o = n1909_o[51];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5694_o = n5693_o;
      7'b0100000: n5694_o = n5693_o;
      7'b0010000: n5694_o = n5693_o;
      7'b0001000: n5694_o = n5692_o;
      7'b0000100: n5694_o = n3858_o;
      7'b0000010: n5694_o = n5693_o;
      7'b0000001: n5694_o = n5693_o;
      default: n5694_o = n5693_o;
    endcase
  assign n5695_o = n3967_o[1];
  assign n5696_o = n1909_o[52];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5697_o = n5696_o;
      7'b0100000: n5697_o = n5696_o;
      7'b0010000: n5697_o = n5696_o;
      7'b0001000: n5697_o = n5695_o;
      7'b0000100: n5697_o = n5696_o;
      7'b0000010: n5697_o = n5696_o;
      7'b0000001: n5697_o = n5696_o;
      default: n5697_o = n5696_o;
    endcase
  assign n5698_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5699_o = n5698_o;
      7'b0100000: n5699_o = n5698_o;
      7'b0010000: n5699_o = n5698_o;
      7'b0001000: n5699_o = n4070_o;
      7'b0000100: n5699_o = n5698_o;
      7'b0000010: n5699_o = n5698_o;
      7'b0000001: n5699_o = n5698_o;
      default: n5699_o = n5698_o;
    endcase
  assign n5700_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5701_o = n5700_o;
      7'b0100000: n5701_o = n5700_o;
      7'b0010000: n5701_o = n4831_o;
      7'b0001000: n5701_o = n5700_o;
      7'b0000100: n5701_o = n3930_o;
      7'b0000010: n5701_o = n3823_o;
      7'b0000001: n5701_o = n3721_o;
      default: n5701_o = n5700_o;
    endcase
  assign n5702_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5703_o = n5604_o;
      7'b0100000: n5703_o = n5702_o;
      7'b0010000: n5703_o = n4833_o;
      7'b0001000: n5703_o = n5702_o;
      7'b0000100: n5703_o = n5702_o;
      7'b0000010: n5703_o = n5702_o;
      7'b0000001: n5703_o = n5702_o;
      default: n5703_o = n5702_o;
    endcase
  assign n5704_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5705_o = n5704_o;
      7'b0100000: n5705_o = n5704_o;
      7'b0010000: n5705_o = n4836_o;
      7'b0001000: n5705_o = n5704_o;
      7'b0000100: n5705_o = n3932_o;
      7'b0000010: n5705_o = n5704_o;
      7'b0000001: n5705_o = n3723_o;
      default: n5705_o = n5704_o;
    endcase
  assign n5706_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5707_o = n5606_o;
      7'b0100000: n5707_o = n5706_o;
      7'b0010000: n5707_o = n5706_o;
      7'b0001000: n5707_o = n5706_o;
      7'b0000100: n5707_o = n5706_o;
      7'b0000010: n5707_o = n5706_o;
      7'b0000001: n5707_o = n5706_o;
      default: n5707_o = n5706_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5708_o = n5059_o;
      7'b0100000: n5708_o = n2178_o;
      7'b0010000: n5708_o = n2178_o;
      7'b0001000: n5708_o = n2178_o;
      7'b0000100: n5708_o = n2178_o;
      7'b0000010: n5708_o = n2178_o;
      7'b0000001: n5708_o = n2178_o;
      default: n5708_o = n2178_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5709_o = n5608_o;
      7'b0100000: n5709_o = n2019_o;
      7'b0010000: n5709_o = n2019_o;
      7'b0001000: n5709_o = n2019_o;
      7'b0000100: n5709_o = n2019_o;
      7'b0000010: n5709_o = n2019_o;
      7'b0000001: n5709_o = n2019_o;
      default: n5709_o = n2019_o;
    endcase
  assign n5710_o = n1909_o[67];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5711_o = n5710_o;
      7'b0100000: n5711_o = n5710_o;
      7'b0010000: n5711_o = n4838_o;
      7'b0001000: n5711_o = n5710_o;
      7'b0000100: n5711_o = n5710_o;
      7'b0000010: n5711_o = n5710_o;
      7'b0000001: n5711_o = n5710_o;
      default: n5711_o = n5710_o;
    endcase
  assign n5712_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5713_o = n5712_o;
      7'b0100000: n5713_o = n5712_o;
      7'b0010000: n5713_o = n4840_o;
      7'b0001000: n5713_o = n5712_o;
      7'b0000100: n5713_o = n5712_o;
      7'b0000010: n5713_o = n5712_o;
      7'b0000001: n5713_o = n5712_o;
      default: n5713_o = n5712_o;
    endcase
  assign n5714_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5715_o = n5714_o;
      7'b0100000: n5715_o = n5714_o;
      7'b0010000: n5715_o = n4841_o;
      7'b0001000: n5715_o = n5714_o;
      7'b0000100: n5715_o = n5714_o;
      7'b0000010: n5715_o = n5714_o;
      7'b0000001: n5715_o = n5714_o;
      default: n5715_o = n5714_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5716_o = n2171_o;
      7'b0100000: n5716_o = n2171_o;
      7'b0010000: n5716_o = n4842_o;
      7'b0001000: n5716_o = n2171_o;
      7'b0000100: n5716_o = n2171_o;
      7'b0000010: n5716_o = n2171_o;
      7'b0000001: n5716_o = n2171_o;
      default: n5716_o = n2171_o;
    endcase
  assign n5717_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5718_o = n5610_o;
      7'b0100000: n5718_o = n5717_o;
      7'b0010000: n5718_o = n5717_o;
      7'b0001000: n5718_o = n5717_o;
      7'b0000100: n5718_o = n5717_o;
      7'b0000010: n5718_o = n5717_o;
      7'b0000001: n5718_o = n5717_o;
      default: n5718_o = n5717_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5720_o = n5613_o;
      7'b0100000: n5720_o = n4971_o;
      7'b0010000: n5720_o = n4844_o;
      7'b0001000: n5720_o = 1'b0;
      7'b0000100: n5720_o = 1'b0;
      7'b0000010: n5720_o = 1'b0;
      7'b0000001: n5720_o = 1'b0;
      default: n5720_o = 1'b0;
    endcase
  assign n5721_o = n3726_o[0];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5723_o = 1'b0;
      7'b0100000: n5723_o = 1'b0;
      7'b0010000: n5723_o = 1'b0;
      7'b0001000: n5723_o = 1'b0;
      7'b0000100: n5723_o = 1'b0;
      7'b0000010: n5723_o = n3825_o;
      7'b0000001: n5723_o = n5721_o;
      default: n5723_o = 1'b0;
    endcase
  assign n5724_o = n3726_o[1];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5726_o = n5615_o;
      7'b0100000: n5726_o = 1'b0;
      7'b0010000: n5726_o = n4846_o;
      7'b0001000: n5726_o = 1'b0;
      7'b0000100: n5726_o = n3934_o;
      7'b0000010: n5726_o = 1'b0;
      7'b0000001: n5726_o = n5724_o;
      default: n5726_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5728_o = 1'b0;
      7'b0100000: n5728_o = 1'b0;
      7'b0010000: n5728_o = 1'b0;
      7'b0001000: n5728_o = 1'b0;
      7'b0000100: n5728_o = 1'b0;
      7'b0000010: n5728_o = n3827_o;
      7'b0000001: n5728_o = 1'b0;
      default: n5728_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5730_o = 1'b0;
      7'b0100000: n5730_o = 1'b0;
      7'b0010000: n5730_o = 1'b0;
      7'b0001000: n5730_o = n4072_o;
      7'b0000100: n5730_o = 1'b0;
      7'b0000010: n5730_o = 1'b0;
      7'b0000001: n5730_o = 1'b0;
      default: n5730_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5732_o = 1'b0;
      7'b0100000: n5732_o = 1'b0;
      7'b0010000: n5732_o = n4848_o;
      7'b0001000: n5732_o = 1'b0;
      7'b0000100: n5732_o = 1'b0;
      7'b0000010: n5732_o = 1'b0;
      7'b0000001: n5732_o = 1'b0;
      default: n5732_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5734_o = 1'b0;
      7'b0100000: n5734_o = 1'b0;
      7'b0010000: n5734_o = n4850_o;
      7'b0001000: n5734_o = 1'b0;
      7'b0000100: n5734_o = 1'b0;
      7'b0000010: n5734_o = 1'b0;
      7'b0000001: n5734_o = 1'b0;
      default: n5734_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5736_o = 1'b0;
      7'b0100000: n5736_o = 1'b0;
      7'b0010000: n5736_o = n4852_o;
      7'b0001000: n5736_o = 1'b0;
      7'b0000100: n5736_o = 1'b0;
      7'b0000010: n5736_o = 1'b0;
      7'b0000001: n5736_o = 1'b0;
      default: n5736_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5738_o = 1'b0;
      7'b0100000: n5738_o = 1'b0;
      7'b0010000: n5738_o = 1'b0;
      7'b0001000: n5738_o = n4074_o;
      7'b0000100: n5738_o = 1'b0;
      7'b0000010: n5738_o = 1'b0;
      7'b0000001: n5738_o = 1'b0;
      default: n5738_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5740_o = 1'b0;
      7'b0100000: n5740_o = 1'b0;
      7'b0010000: n5740_o = n4854_o;
      7'b0001000: n5740_o = 1'b0;
      7'b0000100: n5740_o = 1'b0;
      7'b0000010: n5740_o = 1'b0;
      7'b0000001: n5740_o = n3728_o;
      default: n5740_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5742_o = 1'b0;
      7'b0100000: n5742_o = 1'b0;
      7'b0010000: n5742_o = n4856_o;
      7'b0001000: n5742_o = 1'b0;
      7'b0000100: n5742_o = 1'b0;
      7'b0000010: n5742_o = 1'b0;
      7'b0000001: n5742_o = 1'b0;
      default: n5742_o = 1'b0;
    endcase
  assign n5743_o = n5617_o[1:0];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5745_o = n5743_o;
      7'b0100000: n5745_o = 2'b00;
      7'b0010000: n5745_o = 2'b00;
      7'b0001000: n5745_o = 2'b00;
      7'b0000100: n5745_o = 2'b00;
      7'b0000010: n5745_o = 2'b00;
      7'b0000001: n5745_o = 2'b00;
      default: n5745_o = 2'b00;
    endcase
  assign n5746_o = n5617_o[2];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5748_o = n5746_o;
      7'b0100000: n5748_o = n4973_o;
      7'b0010000: n5748_o = n4857_o;
      7'b0001000: n5748_o = n4076_o;
      7'b0000100: n5748_o = n3936_o;
      7'b0000010: n5748_o = n3829_o;
      7'b0000001: n5748_o = n3730_o;
      default: n5748_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5750_o = 1'b0;
      7'b0100000: n5750_o = 1'b0;
      7'b0010000: n5750_o = n4859_o;
      7'b0001000: n5750_o = 1'b0;
      7'b0000100: n5750_o = 1'b0;
      7'b0000010: n5750_o = 1'b0;
      7'b0000001: n5750_o = 1'b0;
      default: n5750_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5621_o)
      7'b1000000: n5751_o = n5618_o;
      7'b0100000: n5751_o = n2180_o;
      7'b0010000: n5751_o = n4860_o;
      7'b0001000: n5751_o = n2180_o;
      7'b0000100: n5751_o = n2180_o;
      7'b0000010: n5751_o = n2180_o;
      7'b0000001: n5751_o = n2180_o;
      default: n5751_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5752_o = n3356_o ? make_berr : n5622_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5753_o = n3356_o ? n3583_o : n5623_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5754_o = n3356_o ? n3584_o : n5624_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5755_o = n3356_o ? n2148_o : n5625_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5756_o = n3356_o ? n2151_o : n5626_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5758_o = n3356_o ? 1'b0 : n5628_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5759_o = n3356_o ? n2015_o : n5629_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5761_o = n3356_o ? 1'b0 : n5631_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5763_o = n3356_o ? 1'b0 : n5633_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5764_o = n3356_o ? n3586_o : n5635_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5765_o = n3356_o ? n3588_o : n5637_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5766_o = n3356_o ? n3589_o : n5639_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5768_o = n3356_o ? 1'b0 : n5641_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5770_o = n3356_o ? n3591_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5772_o = n3356_o ? 1'b0 : n5643_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5773_o = n3356_o ? n3592_o : n5645_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5774_o = n3356_o ? n1906_o : n5646_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5776_o = n3356_o ? 1'b0 : n5648_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5777_o = n3356_o ? n3593_o : n5649_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5778_o = n3356_o ? n3594_o : n5651_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5780_o = n3356_o ? 1'b0 : n5653_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5782_o = n3356_o ? 1'b0 : n5655_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5784_o = n3356_o ? 1'b0 : n5657_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5785_o = n3356_o ? n3595_o : n5659_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5787_o = n3356_o ? 1'b0 : n5661_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5788_o = n3356_o ? n3596_o : n5663_o;
  assign n5789_o = {n5691_o, n5689_o, n5687_o, n5683_o};
  assign n5790_o = {n5707_o, n5705_o, n5703_o, n5701_o, n5699_o, n5697_o, n5694_o};
  assign n5791_o = {n5711_o, n5709_o, n5708_o};
  assign n5792_o = {n5718_o, n5716_o};
  assign n5793_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5794_o = n3356_o ? n5793_o : n5665_o;
  assign n5795_o = n1909_o[20];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5796_o = n3356_o ? n5795_o : n5667_o;
  assign n5797_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5798_o = n3356_o ? n5797_o : n5669_o;
  assign n5799_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5800_o = n3356_o ? n5799_o : n5671_o;
  assign n5801_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5802_o = n3356_o ? n5801_o : n5673_o;
  assign n5803_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5804_o = n3356_o ? n5803_o : n5675_o;
  assign n5805_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5806_o = n3356_o ? n5805_o : n5677_o;
  assign n5807_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5808_o = n3356_o ? n3598_o : n5807_o;
  assign n5809_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5810_o = n3356_o ? n5809_o : n5679_o;
  assign n5811_o = n5789_o[2:0];
  assign n5812_o = n1909_o[48];
  assign n5813_o = {n5812_o, n2166_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5814_o = n3356_o ? n5813_o : n5811_o;
  assign n5815_o = n5789_o[3];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5816_o = n3356_o ? n3600_o : n5815_o;
  assign n5817_o = n5790_o[4:0];
  assign n5818_o = n1909_o[55:51];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5819_o = n3356_o ? n5818_o : n5817_o;
  assign n5820_o = n5790_o[5];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5821_o = n3356_o ? n3602_o : n5820_o;
  assign n5822_o = n5790_o[9:6];
  assign n5823_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5824_o = n3356_o ? n5823_o : n5822_o;
  assign n5825_o = n1909_o[67];
  assign n5826_o = {n5825_o, n2019_o, n2178_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5827_o = n3356_o ? n5826_o : n5791_o;
  assign n5828_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5829_o = n3356_o ? n5828_o : n5713_o;
  assign n5830_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5831_o = n3356_o ? n5830_o : n5715_o;
  assign n5832_o = n1909_o[74];
  assign n5833_o = {n5832_o, n2171_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5834_o = n3356_o ? n5833_o : n5792_o;
  assign n5835_o = {n5726_o, n5723_o};
  assign n5836_o = {n5730_o, n5728_o};
  assign n5837_o = {n5748_o, n5745_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5838_o = n3356_o ? n3604_o : n5720_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5840_o = n3356_o ? 2'b00 : n5835_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5842_o = n3356_o ? 2'b00 : n5836_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5843_o = n3356_o ? n3606_o : n5732_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5845_o = n3356_o ? 1'b0 : n5734_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5847_o = n3356_o ? 1'b0 : n5736_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5849_o = n3356_o ? 1'b0 : n5738_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5851_o = n3356_o ? 1'b0 : n5740_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5853_o = n3356_o ? 1'b0 : n5742_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5855_o = n3356_o ? n3608_o : 1'b0;
  assign n5856_o = n5837_o[1:0];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5858_o = n3356_o ? 2'b00 : n5856_o;
  assign n5859_o = n5837_o[2];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5860_o = n3356_o ? n3610_o : n5859_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5861_o = n3356_o ? n3612_o : n5750_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5862_o = n3356_o ? n2180_o : n5751_o;
  /* TG68KdotC_Kernel.vhd:1965:25  */
  assign n5864_o = n2185_o == 4'b0100;
  /* TG68KdotC_Kernel.vhd:2644:50  */
  assign n5865_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2644:62  */
  assign n5867_o = n5865_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2645:58  */
  assign n5868_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2645:70  */
  assign n5870_o = n5868_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2646:57  */
  assign n5874_o = decodeopc ? 1'b1 : 1'b0;
  assign n5875_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5876_o = n6071_o ? 1'b1 : n5875_o;
  /* TG68KdotC_Kernel.vhd:2646:57  */
  assign n5878_o = decodeopc ? 7'b0011001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2651:61  */
  assign n5879_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2651:73  */
  assign n5881_o = n5879_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:2651:91  */
  assign n5882_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2651:103  */
  assign n5884_o = n5882_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2651:118  */
  assign n5885_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:2651:130  */
  assign n5887_o = n5885_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2651:109  */
  assign n5888_o = n5884_o | n5887_o;
  /* TG68KdotC_Kernel.vhd:2651:80  */
  assign n5889_o = n5888_o & n5881_o;
  /* TG68KdotC_Kernel.vhd:2652:63  */
  assign n5890_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2653:74  */
  assign n5891_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2653:86  */
  assign n5893_o = n5891_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2655:90  */
  assign n5894_o = opcode[0];
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5896_o = n5975_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2654:73  */
  assign n5897_o = n5894_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5899_o = n5980_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2661:73  */
  assign n5901_o = decodeopc ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2653:65  */
  assign n5902_o = n5893_o ? n2026_o : n5901_o;
  /* TG68KdotC_Kernel.vhd:2653:65  */
  assign n5903_o = n5897_o & n5893_o;
  /* TG68KdotC_Kernel.vhd:2653:65  */
  assign n5904_o = decodeopc & n5893_o;
  /* TG68KdotC_Kernel.vhd:2665:99  */
  assign n5905_o = ~decodeopc;
  /* TG68KdotC_Kernel.vhd:2665:86  */
  assign n5906_o = n5905_o & exe_condition;
  /* TG68KdotC_Kernel.vhd:2665:65  */
  assign n5909_o = n5906_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2665:65  */
  assign n5912_o = n5906_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5913_o = n5966_o ? n5902_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5916_o = n5890_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5918_o = n5890_o ? n5909_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5920_o = n5890_o ? n5912_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5921_o = n5903_o & n5890_o;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5922_o = n5904_o & n5890_o;
  /* TG68KdotC_Kernel.vhd:2673:62  */
  assign n5923_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2673:74  */
  assign n5925_o = n5923_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2673:91  */
  assign n5926_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2673:103  */
  assign n5928_o = n5926_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2673:82  */
  assign n5929_o = n5925_o | n5928_o;
  /* TG68KdotC_Kernel.vhd:2678:63  */
  assign n5931_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2678:80  */
  assign n5933_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2678:71  */
  assign n5934_o = n5933_o & n5931_o;
  /* TG68KdotC_Kernel.vhd:2678:99  */
  assign n5935_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2678:86  */
  assign n5936_o = n5935_o & n5934_o;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5938_o = n5945_o ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2681:66  */
  assign n5939_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2681:78  */
  assign n5941_o = n5939_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2681:57  */
  assign n5944_o = n5941_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5945_o = n5936_o & n5929_o;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5947_o = n5929_o ? 2'b00 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5950_o = n5929_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5953_o = n5929_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5956_o = n5929_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5959_o = n5929_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5961_o = n5929_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5963_o = n5929_o ? n5944_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5964_o = n5889_o ? make_berr : n5938_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5965_o = n5889_o ? n1921_o : n5947_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5966_o = n5890_o & n5889_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5968_o = n5889_o ? 1'b0 : n5950_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5969_o = n5889_o ? n5916_o : n5953_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5971_o = n5889_o ? n5918_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5972_o = n5889_o ? n5920_o : n5956_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5974_o = n5889_o ? 1'b0 : n5959_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5975_o = n5921_o & n5889_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5977_o = n5889_o ? 1'b0 : n5961_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5979_o = n5889_o ? 1'b0 : n5963_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5980_o = n5922_o & n5889_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5981_o = n5870_o ? make_berr : n5964_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5982_o = n5870_o ? n1921_o : n5965_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5983_o = n5870_o ? n2026_o : n5913_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5985_o = n5870_o ? n5874_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5987_o = n5870_o ? 1'b0 : n5968_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5989_o = n5870_o ? 1'b0 : n5969_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5991_o = n5870_o ? 1'b0 : n5971_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5993_o = n5870_o ? 1'b0 : n5972_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5995_o = n5870_o ? 1'b0 : n5974_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5997_o = decodeopc & n5870_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5998_o = n5870_o ? n2171_o : n5896_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n6000_o = n5870_o ? 1'b0 : n5977_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n6002_o = n5870_o ? 1'b0 : n5979_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n6003_o = n5870_o ? n5878_o : n5899_o;
  /* TG68KdotC_Kernel.vhd:2689:58  */
  assign n6004_o = opcode[7:3];
  /* TG68KdotC_Kernel.vhd:2689:70  */
  assign n6006_o = n6004_o != 5'b00001;
  /* TG68KdotC_Kernel.vhd:2690:59  */
  assign n6007_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2690:71  */
  assign n6009_o = n6007_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2690:88  */
  assign n6010_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2690:100  */
  assign n6012_o = n6010_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2690:79  */
  assign n6013_o = n6009_o | n6012_o;
  /* TG68KdotC_Kernel.vhd:2689:80  */
  assign n6014_o = n6013_o & n6006_o;
  /* TG68KdotC_Kernel.vhd:2692:66  */
  assign n6015_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2692:78  */
  assign n6017_o = n6015_o == 3'b001;
  assign n6019_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6020_o = n6047_o ? 1'b1 : n6019_o;
  /* TG68KdotC_Kernel.vhd:2695:66  */
  assign n6021_o = opcode[8];
  assign n6023_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6024_o = n6049_o ? 1'b1 : n6023_o;
  /* TG68KdotC_Kernel.vhd:2702:66  */
  assign n6028_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2702:78  */
  assign n6030_o = n6028_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2702:57  */
  assign n6033_o = n6030_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6036_o = n6014_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6039_o = n6014_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6042_o = n6014_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6045_o = n6014_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6047_o = n6017_o & n6014_o;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6049_o = n6021_o & n6014_o;
  assign n6050_o = {1'b1, 1'b1};
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6052_o = n6014_o ? n6050_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6054_o = n6014_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n6056_o = n6014_o ? n6033_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6057_o = n5867_o ? n5981_o : make_berr;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6058_o = n5867_o ? n5982_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6059_o = n5867_o ? n5983_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6061_o = n5867_o ? n5985_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6062_o = n5867_o ? n5987_o : n6036_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6063_o = n5867_o ? n5989_o : n6039_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6065_o = n5867_o ? n5991_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6066_o = n5867_o ? n5993_o : n6042_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6067_o = n5867_o ? n5995_o : n6045_o;
  assign n6068_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6069_o = n5867_o ? n6068_o : n6020_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6071_o = n5997_o & n5867_o;
  assign n6072_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6073_o = n5867_o ? n6072_o : n6024_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6074_o = n5867_o ? n5998_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6076_o = n5867_o ? 2'b00 : n6052_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6078_o = n5867_o ? n6000_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6080_o = n5867_o ? 1'b0 : n6054_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6081_o = n5867_o ? n6002_o : n6056_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n6082_o = n5867_o ? n6003_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2643:25  */
  assign n6084_o = n2185_o == 4'b0101;
  /* TG68KdotC_Kernel.vhd:2715:47  */
  assign n6086_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2716:50  */
  assign n6087_o = opcode[11:8];
  /* TG68KdotC_Kernel.vhd:2716:63  */
  assign n6089_o = n6087_o == 4'b0001;
  /* TG68KdotC_Kernel.vhd:2719:58  */
  assign n6091_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2719:70  */
  assign n6093_o = n6091_o == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:2722:61  */
  assign n6095_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2722:73  */
  assign n6097_o = n6095_o == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:2722:49  */
  assign n6099_o = n6097_o ? n2026_o : 2'b11;
  /* TG68KdotC_Kernel.vhd:2722:49  */
  assign n6102_o = n6097_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2722:49  */
  assign n6105_o = n6097_o ? 7'b0010111 : 7'b0010110;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n6106_o = n6093_o ? n2026_o : n6099_o;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n6108_o = n6093_o ? 1'b0 : n6102_o;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n6109_o = n6093_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n6111_o = n6093_o ? 7'b0010111 : n6105_o;
  /* TG68KdotC_Kernel.vhd:2730:58  */
  assign n6112_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2730:70  */
  assign n6114_o = n6112_o == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:2733:61  */
  assign n6116_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2733:73  */
  assign n6118_o = n6116_o == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:2733:49  */
  assign n6120_o = n6118_o ? n2026_o : 2'b01;
  /* TG68KdotC_Kernel.vhd:2730:49  */
  assign n6121_o = n6114_o ? n2026_o : n6120_o;
  /* TG68KdotC_Kernel.vhd:2730:49  */
  assign n6122_o = n6114_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n6123_o = n6089_o ? n6106_o : n6121_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n6125_o = n6136_o ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n6127_o = n6089_o ? n6108_o : 1'b0;
  assign n6128_o = n2162_o[1];
  assign n6129_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6130_o = n2037_o ? n6128_o : n6129_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n6131_o = n6089_o ? 1'b1 : n6130_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n6132_o = n6089_o ? n6109_o : n6122_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n6134_o = n6089_o ? n6111_o : 7'b0010101;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n6135_o = n6086_o ? n6123_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n6136_o = n6089_o & n6086_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n6138_o = n6086_o ? n6127_o : 1'b0;
  assign n6139_o = n2162_o[1];
  assign n6140_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6141_o = n2037_o ? n6139_o : n6140_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n6142_o = n6086_o ? n6131_o : n6141_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n6143_o = n6086_o ? n6132_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n6144_o = n6086_o ? n6134_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2712:25  */
  assign n6146_o = n2185_o == 4'b0110;
  /* TG68KdotC_Kernel.vhd:2744:42  */
  assign n6147_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2744:45  */
  assign n6148_o = ~n6147_o;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6153_o = n6148_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6156_o = n6148_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6159_o = n6148_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6162_o = n6148_o ? 1'b0 : 1'b1;
  assign n6163_o = {1'b1, 1'b1};
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6165_o = n6148_o ? n6163_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6167_o = n6148_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2743:25  */
  assign n6169_o = n2185_o == 4'b0111;
  /* TG68KdotC_Kernel.vhd:2757:42  */
  assign n6170_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2757:54  */
  assign n6172_o = n6170_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2759:50  */
  assign n6173_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2759:62  */
  assign n6175_o = n6173_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2758:56  */
  assign n6177_o = n6175_o & 1'b1;
  /* TG68KdotC_Kernel.vhd:2759:81  */
  assign n6178_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2759:93  */
  assign n6180_o = n6178_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2759:111  */
  assign n6181_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2759:123  */
  assign n6183_o = n6181_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2759:102  */
  assign n6184_o = n6180_o | n6183_o;
  /* TG68KdotC_Kernel.vhd:2759:70  */
  assign n6185_o = n6184_o & n6177_o;
  /* TG68KdotC_Kernel.vhd:2760:58  */
  assign n6186_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2760:70  */
  assign n6188_o = n6186_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2760:49  */
  assign n6191_o = n6188_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2763:64  */
  assign n6193_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2763:70  */
  assign n6194_o = nextpass & n6193_o;
  /* TG68KdotC_Kernel.vhd:2763:98  */
  assign n6195_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2763:110  */
  assign n6197_o = n6195_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2763:116  */
  assign n6198_o = decodeopc & n6197_o;
  /* TG68KdotC_Kernel.vhd:2763:88  */
  assign n6199_o = n6194_o | n6198_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6201_o = n6455_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6203_o = n6239_o ? 7'b1010101 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2768:59  */
  assign n6204_o = ~z_error;
  /* TG68KdotC_Kernel.vhd:2768:78  */
  assign n6205_o = ~set_v_flag;
  /* TG68KdotC_Kernel.vhd:2768:64  */
  assign n6206_o = n6205_o & n6204_o;
  /* TG68KdotC_Kernel.vhd:2768:49  */
  assign n6209_o = n6206_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2772:75  */
  assign n6210_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2772:87  */
  assign n6212_o = n6210_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2772:93  */
  assign n6213_o = decodeopc & n6212_o;
  /* TG68KdotC_Kernel.vhd:2772:65  */
  assign n6214_o = nextpass | n6213_o;
  /* TG68KdotC_Kernel.vhd:2772:49  */
  assign n6217_o = n6214_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6219_o = n6185_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6220_o = n6199_o & n6185_o;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6222_o = n6185_o ? n6191_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6225_o = n6185_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6227_o = n6185_o ? n6217_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6230_o = n6185_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6233_o = n6185_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6236_o = n6185_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6238_o = n6185_o ? n6209_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6239_o = n6199_o & n6185_o;
  /* TG68KdotC_Kernel.vhd:2780:45  */
  assign n6240_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2780:63  */
  assign n6241_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2780:75  */
  assign n6243_o = n6241_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2780:53  */
  assign n6244_o = n6243_o & n6240_o;
  /* TG68KdotC_Kernel.vhd:2781:50  */
  assign n6245_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2781:62  */
  assign n6247_o = n6245_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2786:53  */
  assign n6251_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2786:65  */
  assign n6253_o = n6251_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2786:80  */
  assign n6254_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2786:92  */
  assign n6256_o = n6254_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2786:71  */
  assign n6257_o = n6253_o | n6256_o;
  /* TG68KdotC_Kernel.vhd:2790:58  */
  assign n6260_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2790:71  */
  assign n6262_o = n6260_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2790:49  */
  assign n6267_o = n6262_o ? 2'b01 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2790:49  */
  assign n6269_o = n6262_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2790:49  */
  assign n6271_o = n6262_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2797:58  */
  assign n6272_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2797:61  */
  assign n6273_o = ~n6272_o;
  /* TG68KdotC_Kernel.vhd:2798:66  */
  assign n6274_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2798:79  */
  assign n6276_o = n6274_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2798:57  */
  assign n6279_o = n6276_o ? 2'b00 : 2'b01;
  assign n6283_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6284_o = n6325_o ? 1'b1 : n6283_o;
  assign n6285_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6286_o = n6329_o ? 1'b1 : n6285_o;
  /* TG68KdotC_Kernel.vhd:2805:57  */
  assign n6288_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2813:57  */
  assign n6290_o = decodeopc ? 1'b1 : n2154_o;
  /* TG68KdotC_Kernel.vhd:2813:57  */
  assign n6292_o = decodeopc ? 7'b0011110 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6293_o = n6309_o ? n6279_o : datatype;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6296_o = n6273_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6299_o = n6273_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6300_o = n6273_o ? n2154_o : n6290_o;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6302_o = decodeopc & n6273_o;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6304_o = decodeopc & n6273_o;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6306_o = n6273_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6307_o = n6273_o ? n6288_o : n6292_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6308_o = n6257_o ? n6267_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6309_o = n6273_o & n6257_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6311_o = n6257_o ? n6296_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6314_o = n6257_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6316_o = n6257_o ? n6299_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6317_o = n6257_o ? n6300_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6320_o = n6257_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6323_o = n6257_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6325_o = n6302_o & n6257_o;
  assign n6326_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6327_o = n6257_o ? 1'b1 : n6326_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6329_o = n6304_o & n6257_o;
  assign n6330_o = {n6271_o, n6269_o};
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6332_o = n6257_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6334_o = n6257_o ? n6306_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6336_o = n6257_o ? n6330_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6337_o = n6257_o ? n6307_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6338_o = n6247_o ? n1921_o : n6308_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6339_o = n6247_o ? datatype : n6293_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6341_o = n6247_o ? 1'b0 : n6311_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6343_o = n6247_o ? 1'b0 : n6314_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6345_o = n6247_o ? 1'b0 : n6316_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6346_o = n6247_o ? n2154_o : n6317_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6348_o = n6247_o ? 1'b0 : n6320_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6350_o = n6247_o ? 1'b0 : n6323_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6353_o = n6247_o ? 1'b1 : 1'b0;
  assign n6354_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6355_o = n6247_o ? n6354_o : n6284_o;
  assign n6356_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6357_o = n6247_o ? n6356_o : n6327_o;
  assign n6358_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6359_o = n6437_o ? 1'b1 : n6358_o;
  assign n6360_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6361_o = n6247_o ? n6360_o : n6286_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6363_o = n6247_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6365_o = n6247_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6367_o = n6247_o ? 1'b0 : n6332_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6369_o = n6247_o ? 1'b0 : n6334_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6371_o = n6247_o ? 2'b00 : n6336_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6372_o = n6247_o ? n2180_o : n6337_o;
  /* TG68KdotC_Kernel.vhd:2823:50  */
  assign n6373_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2823:62  */
  assign n6375_o = n6373_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:2824:52  */
  assign n6376_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2824:55  */
  assign n6377_o = ~n6376_o;
  /* TG68KdotC_Kernel.vhd:2824:70  */
  assign n6378_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2824:82  */
  assign n6380_o = n6378_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2824:60  */
  assign n6381_o = n6380_o & n6377_o;
  /* TG68KdotC_Kernel.vhd:2824:101  */
  assign n6382_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2824:113  */
  assign n6384_o = n6382_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2824:131  */
  assign n6385_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2824:143  */
  assign n6387_o = n6385_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2824:122  */
  assign n6388_o = n6384_o | n6387_o;
  /* TG68KdotC_Kernel.vhd:2824:90  */
  assign n6389_o = n6388_o & n6381_o;
  /* TG68KdotC_Kernel.vhd:2825:51  */
  assign n6390_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2825:69  */
  assign n6391_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2825:81  */
  assign n6393_o = n6391_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2825:59  */
  assign n6394_o = n6393_o & n6390_o;
  /* TG68KdotC_Kernel.vhd:2825:99  */
  assign n6395_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2825:111  */
  assign n6397_o = n6395_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2825:128  */
  assign n6398_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2825:140  */
  assign n6400_o = n6398_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2825:119  */
  assign n6401_o = n6397_o | n6400_o;
  /* TG68KdotC_Kernel.vhd:2825:88  */
  assign n6402_o = n6401_o & n6394_o;
  /* TG68KdotC_Kernel.vhd:2824:151  */
  assign n6403_o = n6389_o | n6402_o;
  /* TG68KdotC_Kernel.vhd:2823:69  */
  assign n6404_o = n6403_o & n6375_o;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6408_o = n6404_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6411_o = n6404_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6414_o = n6404_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6416_o = n6404_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6417_o = n6244_o ? n6338_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6418_o = n6244_o ? n6339_o : datatype;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6420_o = n6244_o ? n6341_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6422_o = n6244_o ? n6343_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6424_o = n6244_o ? n6345_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6425_o = n6244_o ? n6346_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6426_o = n6244_o ? n6348_o : n6408_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6427_o = n6244_o ? n6350_o : n6411_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6429_o = n6244_o ? 1'b0 : n6414_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6431_o = n6244_o ? n6353_o : 1'b0;
  assign n6432_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6433_o = n6244_o ? n6355_o : n6432_o;
  assign n6434_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6435_o = n6244_o ? n6357_o : n6434_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6437_o = n6247_o & n6244_o;
  assign n6438_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6439_o = n6244_o ? n6361_o : n6438_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6441_o = n6244_o ? n6363_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6443_o = n6244_o ? 1'b0 : n6416_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6445_o = n6244_o ? n6365_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6447_o = n6244_o ? n6367_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6449_o = n6244_o ? n6369_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6451_o = n6244_o ? n6371_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6452_o = n6244_o ? n6372_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6453_o = n6172_o ? n6219_o : n6417_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6454_o = n6172_o ? datatype : n6418_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6455_o = n6220_o & n6172_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6457_o = n6172_o ? n6222_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6459_o = n6172_o ? 1'b0 : n6420_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6460_o = n6172_o ? n6225_o : n6422_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6461_o = n6172_o ? n6227_o : n6424_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6462_o = n6172_o ? n2154_o : n6425_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6463_o = n6172_o ? n6230_o : n6426_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6464_o = n6172_o ? n6233_o : n6427_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6466_o = n6172_o ? n6236_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6468_o = n6172_o ? 1'b0 : n6429_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6470_o = n6172_o ? 1'b0 : n6431_o;
  assign n6471_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6472_o = n6172_o ? n6471_o : n6433_o;
  assign n6473_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6474_o = n6172_o ? n6473_o : n6435_o;
  assign n6475_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6476_o = n6172_o ? n6475_o : n6359_o;
  assign n6477_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6478_o = n6172_o ? n6477_o : n6439_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6480_o = n6172_o ? 1'b0 : n6441_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6482_o = n6172_o ? 1'b0 : n6443_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6484_o = n6172_o ? 1'b0 : n6445_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6486_o = n6172_o ? 1'b0 : n6447_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6487_o = n6172_o ? n6238_o : n6449_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6489_o = n6172_o ? 2'b00 : n6451_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6490_o = n6172_o ? n6203_o : n6452_o;
  /* TG68KdotC_Kernel.vhd:2756:25  */
  assign n6492_o = n2185_o == 4'b1000;
  /* TG68KdotC_Kernel.vhd:2836:42  */
  assign n6493_o = opcode[8:3];
  /* TG68KdotC_Kernel.vhd:2836:54  */
  assign n6495_o = n6493_o != 6'b000001;
  /* TG68KdotC_Kernel.vhd:2837:45  */
  assign n6496_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2837:48  */
  assign n6497_o = ~n6496_o;
  /* TG68KdotC_Kernel.vhd:2837:62  */
  assign n6498_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2837:74  */
  assign n6500_o = n6498_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2837:53  */
  assign n6501_o = n6497_o | n6500_o;
  /* TG68KdotC_Kernel.vhd:2837:92  */
  assign n6502_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2837:104  */
  assign n6504_o = n6502_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2837:122  */
  assign n6505_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2837:134  */
  assign n6507_o = n6505_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2837:113  */
  assign n6508_o = n6504_o | n6507_o;
  /* TG68KdotC_Kernel.vhd:2837:81  */
  assign n6509_o = n6508_o & n6501_o;
  /* TG68KdotC_Kernel.vhd:2838:43  */
  assign n6510_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2838:62  */
  assign n6511_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2838:74  */
  assign n6513_o = n6511_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2838:91  */
  assign n6514_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2838:103  */
  assign n6516_o = n6514_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2838:82  */
  assign n6517_o = n6513_o | n6516_o;
  /* TG68KdotC_Kernel.vhd:2838:51  */
  assign n6518_o = n6517_o & n6510_o;
  /* TG68KdotC_Kernel.vhd:2837:142  */
  assign n6519_o = n6509_o | n6518_o;
  /* TG68KdotC_Kernel.vhd:2836:65  */
  assign n6520_o = n6519_o & n6495_o;
  /* TG68KdotC_Kernel.vhd:2841:50  */
  assign n6522_o = opcode[14];
  /* TG68KdotC_Kernel.vhd:2841:54  */
  assign n6523_o = ~n6522_o;
  assign n6525_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6526_o = n6600_o ? 1'b1 : n6525_o;
  /* TG68KdotC_Kernel.vhd:2844:50  */
  assign n6527_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2844:62  */
  assign n6529_o = n6527_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2845:58  */
  assign n6530_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2845:61  */
  assign n6531_o = ~n6530_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6533_o = n6575_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2850:58  */
  assign n6535_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2850:49  */
  assign n6538_o = n6535_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2854:49  */
  assign n6542_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2854:49  */
  assign n6545_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2859:58  */
  assign n6546_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2859:76  */
  assign n6547_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2859:88  */
  assign n6549_o = n6547_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2859:66  */
  assign n6550_o = n6549_o & n6546_o;
  /* TG68KdotC_Kernel.vhd:2859:49  */
  assign n6553_o = n6550_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2859:49  */
  assign n6556_o = n6550_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6557_o = n6531_o & n6529_o;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6559_o = n6529_o ? n6538_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6562_o = n6529_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6564_o = n6529_o ? n6542_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6566_o = n6529_o ? n6545_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6568_o = n6529_o ? 1'b0 : n6553_o;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6570_o = n6529_o ? 1'b0 : n6556_o;
  assign n6571_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6572_o = n6598_o ? 1'b1 : n6571_o;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6574_o = n6529_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6575_o = n6557_o & n6520_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6577_o = n6520_o ? n6559_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6579_o = n6520_o ? n6562_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6581_o = n6520_o ? n6564_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6583_o = n6520_o ? n6566_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6586_o = n6520_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6589_o = n6520_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6592_o = n6520_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6594_o = n6520_o ? n6568_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6596_o = n6520_o ? n6570_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6598_o = n6529_o & n6520_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6600_o = n6523_o & n6520_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6602_o = n6520_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6604_o = n6520_o ? n6574_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2835:25  */
  assign n6606_o = n2185_o == 4'b1001;
  /* TG68KdotC_Kernel.vhd:2835:36  */
  assign n6608_o = n2185_o == 4'b1101;
  /* TG68KdotC_Kernel.vhd:2835:36  */
  assign n6609_o = n6606_o | n6608_o;
  /* TG68KdotC_Kernel.vhd:2871:25  */
  assign n6611_o = n2185_o == 4'b1010;
  /* TG68KdotC_Kernel.vhd:2876:42  */
  assign n6612_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2876:54  */
  assign n6614_o = n6612_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2877:50  */
  assign n6615_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2877:62  */
  assign n6617_o = n6615_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2877:80  */
  assign n6618_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2877:92  */
  assign n6620_o = n6618_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2877:71  */
  assign n6621_o = n6617_o | n6620_o;
  /* TG68KdotC_Kernel.vhd:2879:58  */
  assign n6622_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2879:61  */
  assign n6623_o = ~n6622_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6626_o = n6790_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2879:49  */
  assign n6628_o = n6623_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2886:66  */
  assign n6630_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2886:57  */
  assign n6633_o = n6630_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6635_o = setexecopc ? n6633_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6638_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6641_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6644_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6646_o = n6623_o & n6621_o;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6648_o = n6621_o ? n6635_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6650_o = n6621_o ? n6638_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6652_o = n6621_o ? n6641_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6654_o = n6621_o ? n6644_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6657_o = n6621_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6660_o = n6621_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6663_o = n6621_o ? 1'b1 : 1'b0;
  assign n6664_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6665_o = n6621_o ? 1'b1 : n6664_o;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6667_o = n6621_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6669_o = n6621_o ? n6628_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2898:50  */
  assign n6670_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2899:58  */
  assign n6671_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2899:70  */
  assign n6673_o = n6671_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2903:74  */
  assign n6675_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:2903:86  */
  assign n6677_o = n6675_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6679_o = n6779_o ? 1'b1 : n2168_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6683_o = n6769_o ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6684_o = n6774_o ? 1'b1 : n2007_o;
  assign n6685_o = n2162_o[0];
  assign n6686_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6687_o = n2037_o ? n6685_o : n6686_o;
  /* TG68KdotC_Kernel.vhd:2902:57  */
  assign n6688_o = decodeopc ? 1'b1 : n6687_o;
  /* TG68KdotC_Kernel.vhd:2902:57  */
  assign n6689_o = n6677_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6691_o = n6789_o ? 7'b0100010 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2914:66  */
  assign n6694_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2914:78  */
  assign n6696_o = n6694_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2914:95  */
  assign n6697_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2914:107  */
  assign n6699_o = n6697_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2914:86  */
  assign n6700_o = n6696_o | n6699_o;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6704_o = n6700_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6707_o = n6700_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6710_o = n6700_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6713_o = n6700_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6715_o = n6700_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6716_o = decodeopc & n6673_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6718_o = n6673_o ? 1'b0 : n6704_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6720_o = n6673_o ? 1'b0 : n6707_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6722_o = n6673_o ? 1'b1 : n6710_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6724_o = n6673_o ? 1'b0 : n6713_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6725_o = decodeopc & n6673_o;
  assign n6726_o = n2162_o[0];
  assign n6727_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6728_o = n2037_o ? n6726_o : n6727_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6729_o = n6673_o ? n6688_o : n6728_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6730_o = n6689_o & n6673_o;
  assign n6731_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6732_o = n6673_o ? 1'b1 : n6731_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6734_o = n6673_o ? 1'b0 : n6715_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6736_o = n6673_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6738_o = n6673_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6739_o = decodeopc & n6673_o;
  /* TG68KdotC_Kernel.vhd:2924:58  */
  assign n6740_o = opcode[8:3];
  /* TG68KdotC_Kernel.vhd:2924:70  */
  assign n6742_o = n6740_o != 6'b000001;
  /* TG68KdotC_Kernel.vhd:2925:59  */
  assign n6743_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2925:71  */
  assign n6745_o = n6743_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2925:89  */
  assign n6746_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2925:101  */
  assign n6748_o = n6746_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2925:80  */
  assign n6749_o = n6745_o | n6748_o;
  /* TG68KdotC_Kernel.vhd:2924:81  */
  assign n6750_o = n6749_o & n6742_o;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6755_o = n6750_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6758_o = n6750_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6761_o = n6750_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6764_o = n6750_o ? 1'b1 : 1'b0;
  assign n6765_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6766_o = n6750_o ? 1'b1 : n6765_o;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6768_o = n6750_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6769_o = n6716_o & n6670_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6770_o = n6670_o ? n6718_o : n6755_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6771_o = n6670_o ? n6720_o : n6758_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6772_o = n6670_o ? n6722_o : n6761_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6773_o = n6670_o ? n6724_o : n6764_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6774_o = n6725_o & n6670_o;
  assign n6775_o = n2162_o[0];
  assign n6776_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6777_o = n2037_o ? n6775_o : n6776_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6778_o = n6670_o ? n6729_o : n6777_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6779_o = n6730_o & n6670_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6780_o = n6670_o ? n6732_o : n6766_o;
  assign n6781_o = {n6736_o, n6734_o};
  assign n6782_o = n6781_o[0];
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6784_o = n6670_o ? n6782_o : 1'b0;
  assign n6785_o = n6781_o[1];
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6786_o = n6670_o ? n6785_o : n6768_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6788_o = n6670_o ? n6738_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6789_o = n6739_o & n6670_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6790_o = n6646_o & n6614_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6791_o = n6614_o ? n2026_o : n6683_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6793_o = n6614_o ? n6648_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6795_o = n6614_o ? n6650_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6797_o = n6614_o ? n6652_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6799_o = n6614_o ? n6654_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6800_o = n6614_o ? n6657_o : n6770_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6801_o = n6614_o ? n6660_o : n6771_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6802_o = n6614_o ? n6663_o : n6772_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6804_o = n6614_o ? 1'b0 : n6773_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6805_o = n6614_o ? n2007_o : n6684_o;
  assign n6806_o = n2162_o[0];
  assign n6807_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6808_o = n2037_o ? n6806_o : n6807_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6809_o = n6614_o ? n6808_o : n6778_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6810_o = n6614_o ? n2168_o : n6679_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6811_o = n6614_o ? n6665_o : n6780_o;
  assign n6812_o = {n6786_o, n6784_o};
  assign n6813_o = n6812_o[0];
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6815_o = n6614_o ? 1'b0 : n6813_o;
  assign n6816_o = n6812_o[1];
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6817_o = n6614_o ? n6667_o : n6816_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6819_o = n6614_o ? n6669_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6821_o = n6614_o ? 1'b0 : n6788_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6822_o = n6614_o ? n2180_o : n6691_o;
  /* TG68KdotC_Kernel.vhd:2875:25  */
  assign n6824_o = n2185_o == 4'b1011;
  /* TG68KdotC_Kernel.vhd:2939:42  */
  assign n6825_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2939:54  */
  assign n6827_o = n6825_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2941:50  */
  assign n6828_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2941:62  */
  assign n6830_o = n6828_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2940:56  */
  assign n6832_o = n6830_o & 1'b1;
  /* TG68KdotC_Kernel.vhd:2941:81  */
  assign n6833_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2941:93  */
  assign n6835_o = n6833_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2941:111  */
  assign n6836_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2941:123  */
  assign n6838_o = n6836_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2941:102  */
  assign n6839_o = n6835_o | n6838_o;
  /* TG68KdotC_Kernel.vhd:2941:70  */
  assign n6840_o = n6839_o & n6832_o;
  /* TG68KdotC_Kernel.vhd:2942:58  */
  assign n6841_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2942:70  */
  assign n6843_o = n6841_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2942:49  */
  assign n6846_o = n6843_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2945:64  */
  assign n6848_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2945:70  */
  assign n6849_o = nextpass & n6848_o;
  /* TG68KdotC_Kernel.vhd:2945:98  */
  assign n6850_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2945:110  */
  assign n6852_o = n6850_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2945:116  */
  assign n6853_o = decodeopc & n6852_o;
  /* TG68KdotC_Kernel.vhd:2945:88  */
  assign n6854_o = n6849_o | n6853_o;
  /* TG68KdotC_Kernel.vhd:2945:49  */
  assign n6858_o = n6854_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2945:49  */
  assign n6860_o = n6854_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2958:77  */
  assign n6862_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2958:89  */
  assign n6864_o = n6862_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2958:95  */
  assign n6865_o = decodeopc & n6864_o;
  /* TG68KdotC_Kernel.vhd:2958:67  */
  assign n6866_o = nextpass | n6865_o;
  /* TG68KdotC_Kernel.vhd:2958:49  */
  assign n6869_o = n6866_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6872_o = setexecopc ? 2'b10 : 2'b01;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6874_o = n6840_o ? n6872_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6876_o = n6840_o ? n6846_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6879_o = n6840_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6881_o = n6840_o ? n6869_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6884_o = n6840_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6887_o = n6840_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6890_o = n6840_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6892_o = n6840_o ? n6858_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6894_o = n6840_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6896_o = n6840_o ? n6860_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:45  */
  assign n6897_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2969:63  */
  assign n6898_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2969:75  */
  assign n6900_o = n6898_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2969:53  */
  assign n6901_o = n6900_o & n6897_o;
  /* TG68KdotC_Kernel.vhd:2970:50  */
  assign n6902_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2970:62  */
  assign n6904_o = n6902_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2975:58  */
  assign n6907_o = opcode[7:4];
  /* TG68KdotC_Kernel.vhd:2975:70  */
  assign n6909_o = n6907_o == 4'b0100;
  /* TG68KdotC_Kernel.vhd:2975:87  */
  assign n6910_o = opcode[7:3];
  /* TG68KdotC_Kernel.vhd:2975:99  */
  assign n6912_o = n6910_o == 5'b10001;
  /* TG68KdotC_Kernel.vhd:2975:78  */
  assign n6913_o = n6909_o | n6912_o;
  /* TG68KdotC_Kernel.vhd:2980:66  */
  assign n6917_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2980:84  */
  assign n6918_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2980:74  */
  assign n6919_o = n6918_o & n6917_o;
  /* TG68KdotC_Kernel.vhd:2980:57  */
  assign n6922_o = n6919_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2980:57  */
  assign n6925_o = n6919_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6927_o = n6933_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2984:57  */
  assign n6930_o = decodeopc ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6932_o = n6913_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6933_o = decodeopc & n6913_o;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6935_o = n6913_o ? n6922_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6937_o = n6913_o ? n6925_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6939_o = n6913_o ? n6930_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6942_o = n6913_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6945_o = n6913_o ? 1'b0 : 1'b1;
  assign n6946_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6947_o = n6913_o ? 1'b1 : n6946_o;
  assign n6948_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6949_o = n6913_o ? 1'b1 : n6948_o;
  assign n6950_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6951_o = n6913_o ? 1'b1 : n6950_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6952_o = n6904_o ? n1921_o : n6932_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6953_o = n6904_o ? n2026_o : n6927_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6955_o = n6904_o ? 1'b0 : n6935_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6957_o = n6904_o ? 1'b0 : n6937_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6959_o = n6904_o ? 1'b0 : n6939_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6961_o = n6904_o ? 1'b0 : n6942_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6963_o = n6904_o ? 1'b0 : n6945_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6966_o = n6904_o ? 1'b1 : 1'b0;
  assign n6967_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6968_o = n6904_o ? n6967_o : n6947_o;
  assign n6969_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6970_o = n6904_o ? n6969_o : n6949_o;
  assign n6971_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6972_o = n6904_o ? n6971_o : n6951_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6974_o = n6904_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6976_o = n6904_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:50  */
  assign n6977_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2995:62  */
  assign n6979_o = n6977_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:2996:52  */
  assign n6980_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2996:55  */
  assign n6981_o = ~n6980_o;
  /* TG68KdotC_Kernel.vhd:2996:70  */
  assign n6982_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2996:82  */
  assign n6984_o = n6982_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2996:60  */
  assign n6985_o = n6984_o & n6981_o;
  /* TG68KdotC_Kernel.vhd:2996:101  */
  assign n6986_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2996:113  */
  assign n6988_o = n6986_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2996:131  */
  assign n6989_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2996:143  */
  assign n6991_o = n6989_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2996:122  */
  assign n6992_o = n6988_o | n6991_o;
  /* TG68KdotC_Kernel.vhd:2996:90  */
  assign n6993_o = n6992_o & n6985_o;
  /* TG68KdotC_Kernel.vhd:2997:51  */
  assign n6994_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2997:69  */
  assign n6995_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2997:81  */
  assign n6997_o = n6995_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2997:59  */
  assign n6998_o = n6997_o & n6994_o;
  /* TG68KdotC_Kernel.vhd:2997:99  */
  assign n6999_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2997:111  */
  assign n7001_o = n6999_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2997:128  */
  assign n7002_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2997:140  */
  assign n7004_o = n7002_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2997:119  */
  assign n7005_o = n7001_o | n7004_o;
  /* TG68KdotC_Kernel.vhd:2997:88  */
  assign n7006_o = n7005_o & n6998_o;
  /* TG68KdotC_Kernel.vhd:2996:151  */
  assign n7007_o = n6993_o | n7006_o;
  /* TG68KdotC_Kernel.vhd:2995:69  */
  assign n7008_o = n7007_o & n6979_o;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n7012_o = n7008_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n7015_o = n7008_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n7018_o = n7008_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n7020_o = n7008_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7021_o = n6901_o ? n6952_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7022_o = n6901_o ? n6953_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7024_o = n6901_o ? n6955_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7026_o = n6901_o ? n6957_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7028_o = n6901_o ? n6959_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7029_o = n6901_o ? n6961_o : n7012_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7030_o = n6901_o ? n6963_o : n7015_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7032_o = n6901_o ? 1'b0 : n7018_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7034_o = n6901_o ? n6966_o : 1'b0;
  assign n7035_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7036_o = n6901_o ? n6968_o : n7035_o;
  assign n7037_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7038_o = n6901_o ? n6970_o : n7037_o;
  assign n7039_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7040_o = n6901_o ? n6972_o : n7039_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7042_o = n6901_o ? n6974_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7044_o = n6901_o ? 1'b0 : n7020_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n7046_o = n6901_o ? n6976_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7047_o = n6827_o ? n6874_o : n7021_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7048_o = n6827_o ? n2026_o : n7022_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7050_o = n6827_o ? n6876_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7052_o = n6827_o ? 1'b0 : n7024_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7054_o = n6827_o ? n6879_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7056_o = n6827_o ? 1'b0 : n7026_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7057_o = n6827_o ? n6881_o : n7028_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7058_o = n6827_o ? n6884_o : n7029_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7059_o = n6827_o ? n6887_o : n7030_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7061_o = n6827_o ? n6890_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7063_o = n6827_o ? 1'b0 : n7032_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7065_o = n6827_o ? 1'b0 : n7034_o;
  assign n7066_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7067_o = n6827_o ? n7066_o : n7036_o;
  assign n7068_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7069_o = n6827_o ? n7068_o : n7038_o;
  assign n7070_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7071_o = n6827_o ? n7070_o : n7040_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7073_o = n6827_o ? 1'b0 : n7042_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7075_o = n6827_o ? 1'b0 : n7044_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7077_o = n6827_o ? 1'b0 : n7046_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7079_o = n6827_o ? n6892_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7081_o = n6827_o ? n6894_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n7083_o = n6827_o ? n6896_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2938:25  */
  assign n7085_o = n2185_o == 4'b1100;
  /* TG68KdotC_Kernel.vhd:3008:42  */
  assign n7086_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:3008:54  */
  assign n7088_o = n7086_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:3009:50  */
  assign n7089_o = opcode[11];
  /* TG68KdotC_Kernel.vhd:3009:54  */
  assign n7090_o = ~n7089_o;
  /* TG68KdotC_Kernel.vhd:3010:54  */
  assign n7091_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3010:66  */
  assign n7093_o = n7091_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3010:84  */
  assign n7094_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3010:96  */
  assign n7096_o = n7094_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:3010:113  */
  assign n7097_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3010:125  */
  assign n7099_o = n7097_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3010:104  */
  assign n7100_o = n7096_o | n7099_o;
  /* TG68KdotC_Kernel.vhd:3010:73  */
  assign n7101_o = n7100_o & n7093_o;
  /* TG68KdotC_Kernel.vhd:3018:79  */
  assign n7103_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7106_o = n7391_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n7109_o = n7101_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7110_o = n7408_o ? n7103_o : n1900_o;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n7113_o = n7101_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n7116_o = n7101_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n7119_o = n7101_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n7121_o = n7101_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n7123_o = n7101_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3026:70  */
  assign n7124_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3026:73  */
  assign n7125_o = ~n7124_o;
  /* TG68KdotC_Kernel.vhd:3026:78  */
  assign n7127_o = 1'b1 & n7125_o;
  /* TG68KdotC_Kernel.vhd:3026:63  */
  assign n7129_o = 1'b0 | n7127_o;
  /* TG68KdotC_Kernel.vhd:3027:60  */
  assign n7130_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3027:73  */
  assign n7132_o = n7130_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:3027:88  */
  assign n7133_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3027:101  */
  assign n7135_o = n7133_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:3027:79  */
  assign n7136_o = n7132_o | n7135_o;
  /* TG68KdotC_Kernel.vhd:3027:117  */
  assign n7137_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3027:130  */
  assign n7139_o = n7137_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3027:108  */
  assign n7140_o = n7136_o | n7139_o;
  /* TG68KdotC_Kernel.vhd:3028:59  */
  assign n7141_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:71  */
  assign n7143_o = n7141_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3028:87  */
  assign n7144_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:99  */
  assign n7146_o = n7144_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3028:78  */
  assign n7147_o = n7143_o | n7146_o;
  /* TG68KdotC_Kernel.vhd:3028:115  */
  assign n7148_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:127  */
  assign n7150_o = n7148_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3028:106  */
  assign n7151_o = n7147_o | n7150_o;
  /* TG68KdotC_Kernel.vhd:3028:144  */
  assign n7152_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:156  */
  assign n7154_o = n7152_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3028:173  */
  assign n7155_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3028:185  */
  assign n7157_o = n7155_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3028:163  */
  assign n7158_o = n7157_o & n7154_o;
  /* TG68KdotC_Kernel.vhd:3028:134  */
  assign n7159_o = n7151_o | n7158_o;
  /* TG68KdotC_Kernel.vhd:3027:138  */
  assign n7160_o = n7159_o & n7140_o;
  /* TG68KdotC_Kernel.vhd:3026:94  */
  assign n7161_o = n7129_o | n7160_o;
  /* TG68KdotC_Kernel.vhd:3029:60  */
  assign n7162_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3029:73  */
  assign n7164_o = n7162_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3029:88  */
  assign n7165_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3029:101  */
  assign n7167_o = n7165_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3029:79  */
  assign n7168_o = n7164_o | n7167_o;
  /* TG68KdotC_Kernel.vhd:3029:117  */
  assign n7169_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3029:130  */
  assign n7171_o = n7169_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3029:108  */
  assign n7172_o = n7168_o | n7171_o;
  /* TG68KdotC_Kernel.vhd:3030:59  */
  assign n7173_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3030:71  */
  assign n7175_o = n7173_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3030:87  */
  assign n7176_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3030:99  */
  assign n7178_o = n7176_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3030:78  */
  assign n7179_o = n7175_o | n7178_o;
  /* TG68KdotC_Kernel.vhd:3030:115  */
  assign n7180_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3030:127  */
  assign n7182_o = n7180_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3030:106  */
  assign n7183_o = n7179_o | n7182_o;
  /* TG68KdotC_Kernel.vhd:3030:143  */
  assign n7184_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:3030:155  */
  assign n7186_o = n7184_o == 4'b1111;
  /* TG68KdotC_Kernel.vhd:3030:134  */
  assign n7187_o = n7183_o | n7186_o;
  /* TG68KdotC_Kernel.vhd:3029:138  */
  assign n7188_o = n7187_o & n7172_o;
  /* TG68KdotC_Kernel.vhd:3028:195  */
  assign n7189_o = n7161_o | n7188_o;
  assign n7192_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3034:57  */
  assign n7193_o = decodeopc ? 1'b1 : n7192_o;
  assign n7194_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3034:57  */
  assign n7195_o = decodeopc ? 1'b1 : n7194_o;
  /* TG68KdotC_Kernel.vhd:3034:57  */
  assign n7197_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:3041:66  */
  assign n7199_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:3041:84  */
  assign n7200_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:3041:87  */
  assign n7201_o = ~n7200_o;
  /* TG68KdotC_Kernel.vhd:3041:75  */
  assign n7202_o = n7199_o | n7201_o;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7205_o = n7202_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3044:66  */
  assign n7206_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3044:79  */
  assign n7208_o = n7206_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3044:57  */
  assign n7211_o = n7208_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3047:66  */
  assign n7212_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:79  */
  assign n7214_o = n7212_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:3047:95  */
  assign n7215_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:108  */
  assign n7217_o = n7215_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3047:86  */
  assign n7218_o = n7214_o | n7217_o;
  /* TG68KdotC_Kernel.vhd:3047:124  */
  assign n7219_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:137  */
  assign n7221_o = n7219_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:3047:115  */
  assign n7222_o = n7218_o | n7221_o;
  /* TG68KdotC_Kernel.vhd:3047:153  */
  assign n7223_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:166  */
  assign n7225_o = n7223_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3047:144  */
  assign n7226_o = n7222_o | n7225_o;
  /* TG68KdotC_Kernel.vhd:3047:57  */
  assign n7229_o = n7226_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3051:66  */
  assign n7230_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3051:79  */
  assign n7232_o = n7230_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3051:95  */
  assign n7233_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3051:108  */
  assign n7235_o = n7233_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3051:86  */
  assign n7236_o = n7232_o | n7235_o;
  /* TG68KdotC_Kernel.vhd:3051:124  */
  assign n7237_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3051:137  */
  assign n7239_o = n7237_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3051:115  */
  assign n7240_o = n7236_o | n7239_o;
  /* TG68KdotC_Kernel.vhd:3051:57  */
  assign n7243_o = n7240_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3054:66  */
  assign n7244_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:3054:78  */
  assign n7246_o = n7244_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3055:74  */
  assign n7247_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3055:87  */
  assign n7249_o = n7247_o != 3'b000;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7251_o = n7271_o ? 1'b1 : n7243_o;
  /* TG68KdotC_Kernel.vhd:3058:72  */
  assign n7252_o = exec[42];
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7255_o = n7264_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:3058:65  */
  assign n7258_o = n7252_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3058:65  */
  assign n7261_o = n7252_o ? 1'b1 : 1'b0;
  assign n7262_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7263_o = n7270_o ? 1'b1 : n7262_o;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7264_o = n7252_o & n7246_o;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7266_o = n7246_o ? n7258_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7268_o = n7246_o ? n7261_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7270_o = n7252_o & n7246_o;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7271_o = n7249_o & n7246_o;
  /* TG68KdotC_Kernel.vhd:3065:63  */
  assign n7272_o = set[62];
  /* TG68KdotC_Kernel.vhd:3065:57  */
  assign n7274_o = n7272_o ? 2'b01 : n7255_o;
  /* TG68KdotC_Kernel.vhd:3068:64  */
  assign n7275_o = exec[62];
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7279_o = n7275_o ? 2'b01 : n7274_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7281_o = n7275_o ? 1'b1 : n7266_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7283_o = n7275_o ? 1'b1 : n7268_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7284_o = n7275_o ? 1'b1 : n7263_o;
  assign n7285_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7286_o = n7275_o ? 1'b1 : n7285_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7288_o = n7275_o ? 7'b1010000 : n7197_o;
  /* TG68KdotC_Kernel.vhd:3077:74  */
  assign n7289_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3077:87  */
  assign n7291_o = n7289_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3077:65  */
  assign n7294_o = n7291_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3077:65  */
  assign n7297_o = n7291_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3082:74  */
  assign n7298_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3082:87  */
  assign n7300_o = n7298_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3082:103  */
  assign n7301_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3082:116  */
  assign n7303_o = n7301_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3082:94  */
  assign n7304_o = n7300_o | n7303_o;
  /* TG68KdotC_Kernel.vhd:3082:132  */
  assign n7305_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3082:145  */
  assign n7307_o = n7305_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3082:123  */
  assign n7308_o = n7304_o | n7307_o;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7310_o = n7315_o ? 1'b1 : n7283_o;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7312_o = setexecopc ? n7294_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7314_o = setexecopc ? n7297_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7315_o = n7308_o & setexecopc;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7316_o = n7189_o ? n2026_o : n7279_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7318_o = n7189_o ? 1'b0 : n7229_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7321_o = n7189_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7323_o = n7189_o ? 1'b0 : n7312_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7325_o = n7189_o ? 1'b0 : n7314_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7327_o = n7189_o ? 1'b0 : n7281_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7329_o = n7189_o ? 1'b0 : n7310_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7332_o = n7189_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7335_o = n7189_o ? 1'b1 : 1'b0;
  assign n7336_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7337_o = n7189_o ? n7336_o : n7284_o;
  assign n7338_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7339_o = n7189_o ? n7338_o : n7193_o;
  assign n7340_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7341_o = n7189_o ? n7340_o : n7286_o;
  assign n7342_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7343_o = n7189_o ? n7342_o : n7195_o;
  assign n7344_o = {n7205_o, 1'b1};
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7346_o = n7189_o ? 1'b0 : n7211_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7348_o = n7189_o ? 1'b0 : n7251_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7350_o = n7189_o ? 2'b00 : n7344_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7351_o = n7189_o ? n2180_o : n7288_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7352_o = n7101_o & n7090_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7353_o = n7090_o ? n2026_o : n7316_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7354_o = n7090_o ? n7109_o : n7318_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7356_o = n7090_o ? 1'b0 : n7321_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7358_o = n7090_o ? 1'b0 : n7323_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7360_o = n7090_o ? 1'b0 : n7325_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7362_o = n7090_o ? 1'b0 : n7327_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7364_o = n7090_o ? 1'b0 : n7329_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7365_o = n7101_o & n7090_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7366_o = n7090_o ? n7113_o : n7332_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7367_o = n7090_o ? n7116_o : n7335_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7369_o = n7090_o ? n7119_o : 1'b0;
  assign n7370_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7371_o = n7090_o ? n7370_o : n7337_o;
  assign n7372_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7373_o = n7090_o ? n7372_o : n7339_o;
  assign n7374_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7375_o = n7090_o ? n7374_o : n7341_o;
  assign n7376_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7377_o = n7090_o ? n7376_o : n7343_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7378_o = n7090_o ? n7121_o : n7346_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7380_o = n7090_o ? 1'b0 : n7348_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7382_o = n7090_o ? 2'b00 : n7350_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7384_o = n7090_o ? n7123_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7385_o = n7090_o ? n2180_o : n7351_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7391_o = n7352_o & n7088_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7392_o = n7088_o ? n7353_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7395_o = n7088_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7397_o = n7088_o ? n7354_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7399_o = n7088_o ? n7356_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7401_o = n7088_o ? n7358_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7403_o = n7088_o ? n7360_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7405_o = n7088_o ? n7362_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7407_o = n7088_o ? n7364_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7408_o = n7365_o & n7088_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7410_o = n7088_o ? n7366_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7412_o = n7088_o ? n7367_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7414_o = n7088_o ? n7369_o : 1'b0;
  assign n7415_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7416_o = n7088_o ? n7371_o : n7415_o;
  assign n7417_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7418_o = n7088_o ? n7373_o : n7417_o;
  assign n7419_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7420_o = n7088_o ? n7375_o : n7419_o;
  assign n7421_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7422_o = n7088_o ? n7377_o : n7421_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7424_o = n7088_o ? n7378_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7425_o = n7088_o ? n7380_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7427_o = n7088_o ? n7382_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7428_o = n7088_o ? n7384_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7429_o = n7088_o ? n7385_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:3007:25  */
  assign n7431_o = n2185_o == 4'b1110;
  /* TG68KdotC_Kernel.vhd:3117:39  */
  assign n7432_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3117:57  */
  assign n7433_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:3117:69  */
  assign n7435_o = n7433_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3117:47  */
  assign n7436_o = n7435_o & n7432_o;
  /* TG68KdotC_Kernel.vhd:3118:50  */
  assign n7437_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3118:62  */
  assign n7439_o = n7437_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3118:79  */
  assign n7440_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3118:91  */
  assign n7442_o = n7440_o != 3'b011;
  /* TG68KdotC_Kernel.vhd:3118:69  */
  assign n7443_o = n7442_o & n7439_o;
  /* TG68KdotC_Kernel.vhd:3119:51  */
  assign n7444_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3119:63  */
  assign n7446_o = n7444_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:3119:80  */
  assign n7447_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3119:92  */
  assign n7449_o = n7447_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3119:71  */
  assign n7450_o = n7446_o | n7449_o;
  /* TG68KdotC_Kernel.vhd:3118:99  */
  assign n7451_o = n7450_o & n7443_o;
  /* TG68KdotC_Kernel.vhd:3120:58  */
  assign n7452_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3120:71  */
  assign n7454_o = n7452_o != 3'b000;
  /* TG68KdotC_Kernel.vhd:3122:74  */
  assign n7455_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:3122:77  */
  assign n7456_o = ~n7455_o;
  /* TG68KdotC_Kernel.vhd:3122:92  */
  assign n7457_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3122:104  */
  assign n7459_o = n7457_o != 2'b01;
  /* TG68KdotC_Kernel.vhd:3122:82  */
  assign n7460_o = n7459_o & n7456_o;
  /* TG68KdotC_Kernel.vhd:3122:65  */
  assign n7463_o = n7460_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3122:65  */
  assign n7466_o = n7460_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3121:57  */
  assign n7468_o = svmode ? n7463_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3121:57  */
  assign n7471_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3121:57  */
  assign n7473_o = svmode ? n7466_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3136:57  */
  assign n7476_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3136:57  */
  assign n7479_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3120:49  */
  assign n7481_o = n7454_o ? n7468_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3120:49  */
  assign n7482_o = n7454_o ? n7471_o : n7476_o;
  /* TG68KdotC_Kernel.vhd:3120:49  */
  assign n7483_o = n7454_o ? n7473_o : n7479_o;
  /* TG68KdotC_Kernel.vhd:3118:41  */
  assign n7485_o = n7451_o ? n7481_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3118:41  */
  assign n7487_o = n7451_o ? n7482_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3118:41  */
  assign n7489_o = n7451_o ? n7483_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3148:42  */
  assign n7490_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3148:60  */
  assign n7491_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:3148:72  */
  assign n7493_o = n7491_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3148:50  */
  assign n7494_o = n7493_o & n7490_o;
  /* TG68KdotC_Kernel.vhd:3149:50  */
  assign n7495_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3149:62  */
  assign n7497_o = n7495_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3149:79  */
  assign n7498_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3149:91  */
  assign n7500_o = n7498_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:3149:69  */
  assign n7501_o = n7500_o & n7497_o;
  /* TG68KdotC_Kernel.vhd:3150:51  */
  assign n7502_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3150:63  */
  assign n7504_o = n7502_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:3150:81  */
  assign n7505_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3150:93  */
  assign n7507_o = n7505_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:3151:50  */
  assign n7508_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:3151:62  */
  assign n7510_o = n7508_o != 3'b101;
  /* TG68KdotC_Kernel.vhd:3150:100  */
  assign n7511_o = n7510_o & n7507_o;
  /* TG68KdotC_Kernel.vhd:3150:71  */
  assign n7512_o = n7504_o | n7511_o;
  /* TG68KdotC_Kernel.vhd:3149:99  */
  assign n7513_o = n7512_o & n7501_o;
  /* TG68KdotC_Kernel.vhd:3152:58  */
  assign n7514_o = opcode[5:1];
  /* TG68KdotC_Kernel.vhd:3152:70  */
  assign n7516_o = n7514_o != 5'b11110;
  /* TG68KdotC_Kernel.vhd:3153:66  */
  assign n7517_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3153:79  */
  assign n7519_o = n7517_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3153:95  */
  assign n7520_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3153:108  */
  assign n7522_o = n7520_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:3153:86  */
  assign n7523_o = n7519_o | n7522_o;
  /* TG68KdotC_Kernel.vhd:3155:82  */
  assign n7524_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3155:94  */
  assign n7526_o = n7524_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3155:73  */
  assign n7529_o = n7526_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3155:73  */
  assign n7532_o = n7526_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3154:65  */
  assign n7534_o = svmode ? n7529_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3154:65  */
  assign n7537_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3154:65  */
  assign n7539_o = svmode ? n7532_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3168:65  */
  assign n7542_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3168:65  */
  assign n7545_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3153:57  */
  assign n7547_o = n7523_o ? n7534_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3153:57  */
  assign n7548_o = n7523_o ? n7537_o : n7542_o;
  /* TG68KdotC_Kernel.vhd:3153:57  */
  assign n7549_o = n7523_o ? n7539_o : n7545_o;
  /* TG68KdotC_Kernel.vhd:3152:49  */
  assign n7551_o = n7516_o ? n7547_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3152:49  */
  assign n7553_o = n7516_o ? n7548_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3152:49  */
  assign n7555_o = n7516_o ? n7549_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3149:41  */
  assign n7557_o = n7513_o ? n7551_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3149:41  */
  assign n7559_o = n7513_o ? n7553_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3149:41  */
  assign n7561_o = n7513_o ? n7555_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3148:33  */
  assign n7563_o = n7494_o ? n7557_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3148:33  */
  assign n7565_o = n7494_o ? n7559_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3148:33  */
  assign n7567_o = n7494_o ? n7561_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3117:33  */
  assign n7568_o = n7436_o ? n7485_o : n7563_o;
  /* TG68KdotC_Kernel.vhd:3117:33  */
  assign n7569_o = n7436_o ? n7487_o : n7565_o;
  /* TG68KdotC_Kernel.vhd:3117:33  */
  assign n7570_o = n7436_o ? n7489_o : n7567_o;
  /* TG68KdotC_Kernel.vhd:3116:25  */
  assign n7572_o = n2185_o == 4'b1111;
  assign n7573_o = {n7572_o, n7431_o, n7085_o, n6824_o, n6611_o, n6609_o, n6492_o, n6169_o, n6146_o, n6084_o, n5864_o, n3355_o, n3141_o};
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7574_o = make_berr;
      13'b0100000000000: n7574_o = make_berr;
      13'b0010000000000: n7574_o = make_berr;
      13'b0001000000000: n7574_o = make_berr;
      13'b0000100000000: n7574_o = make_berr;
      13'b0000010000000: n7574_o = make_berr;
      13'b0000001000000: n7574_o = make_berr;
      13'b0000000100000: n7574_o = make_berr;
      13'b0000000010000: n7574_o = make_berr;
      13'b0000000001000: n7574_o = n6057_o;
      13'b0000000000100: n7574_o = n5752_o;
      13'b0000000000010: n7574_o = make_berr;
      13'b0000000000001: n7574_o = make_berr;
      default: n7574_o = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7576_o = n1921_o;
      13'b0100000000000: n7576_o = n7106_o;
      13'b0010000000000: n7576_o = n7047_o;
      13'b0001000000000: n7576_o = n6626_o;
      13'b0000100000000: n7576_o = n1921_o;
      13'b0000010000000: n7576_o = n6533_o;
      13'b0000001000000: n7576_o = n6453_o;
      13'b0000000100000: n7576_o = n6153_o;
      13'b0000000010000: n7576_o = 2'b10;
      13'b0000000001000: n7576_o = n6058_o;
      13'b0000000000100: n7576_o = n5753_o;
      13'b0000000000010: n7576_o = n3314_o;
      13'b0000000000001: n7576_o = n3080_o;
      default: n7576_o = n1921_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7577_o = datatype;
      13'b0100000000000: n7577_o = datatype;
      13'b0010000000000: n7577_o = datatype;
      13'b0001000000000: n7577_o = datatype;
      13'b0000100000000: n7577_o = datatype;
      13'b0000010000000: n7577_o = datatype;
      13'b0000001000000: n7577_o = n6454_o;
      13'b0000000100000: n7577_o = datatype;
      13'b0000000010000: n7577_o = datatype;
      13'b0000000001000: n7577_o = datatype;
      13'b0000000000100: n7577_o = datatype;
      13'b0000000000010: n7577_o = datatype;
      13'b0000000000001: n7577_o = datatype;
      default: n7577_o = datatype;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7578_o = n2026_o;
      13'b0100000000000: n7578_o = n7392_o;
      13'b0010000000000: n7578_o = n7048_o;
      13'b0001000000000: n7578_o = n6791_o;
      13'b0000100000000: n7578_o = n2026_o;
      13'b0000010000000: n7578_o = n2026_o;
      13'b0000001000000: n7578_o = n6201_o;
      13'b0000000100000: n7578_o = n2026_o;
      13'b0000000010000: n7578_o = n6135_o;
      13'b0000000001000: n7578_o = n6059_o;
      13'b0000000000100: n7578_o = n5754_o;
      13'b0000000000010: n7578_o = n3304_o;
      13'b0000000000001: n7578_o = n3081_o;
      default: n7578_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7579_o = n2148_o;
      13'b0100000000000: n7579_o = n2148_o;
      13'b0010000000000: n7579_o = n2148_o;
      13'b0001000000000: n7579_o = n2148_o;
      13'b0000100000000: n7579_o = n2148_o;
      13'b0000010000000: n7579_o = n2148_o;
      13'b0000001000000: n7579_o = n2148_o;
      13'b0000000100000: n7579_o = n2148_o;
      13'b0000000010000: n7579_o = n2148_o;
      13'b0000000001000: n7579_o = n2148_o;
      13'b0000000000100: n7579_o = n5755_o;
      13'b0000000000010: n7579_o = n2148_o;
      13'b0000000000001: n7579_o = n2148_o;
      default: n7579_o = n2148_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7581_o = 1'b0;
      13'b0100000000000: n7581_o = 1'b0;
      13'b0010000000000: n7581_o = n7050_o;
      13'b0001000000000: n7581_o = 1'b0;
      13'b0000100000000: n7581_o = 1'b0;
      13'b0000010000000: n7581_o = 1'b0;
      13'b0000001000000: n7581_o = n6457_o;
      13'b0000000100000: n7581_o = 1'b0;
      13'b0000000010000: n7581_o = 1'b0;
      13'b0000000001000: n7581_o = 1'b0;
      13'b0000000000100: n7581_o = 1'b0;
      13'b0000000000010: n7581_o = 1'b0;
      13'b0000000000001: n7581_o = 1'b0;
      default: n7581_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7582_o = n2151_o;
      13'b0100000000000: n7582_o = n2151_o;
      13'b0010000000000: n7582_o = n2151_o;
      13'b0001000000000: n7582_o = n2151_o;
      13'b0000100000000: n7582_o = n2151_o;
      13'b0000010000000: n7582_o = n2151_o;
      13'b0000001000000: n7582_o = n2151_o;
      13'b0000000100000: n7582_o = n2151_o;
      13'b0000000010000: n7582_o = n2151_o;
      13'b0000000001000: n7582_o = n2151_o;
      13'b0000000000100: n7582_o = n5756_o;
      13'b0000000000010: n7582_o = n3305_o;
      13'b0000000000001: n7582_o = n2151_o;
      default: n7582_o = n2151_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7584_o = 1'b0;
      13'b0100000000000: n7584_o = n7395_o;
      13'b0010000000000: n7584_o = 1'b0;
      13'b0001000000000: n7584_o = 1'b0;
      13'b0000100000000: n7584_o = 1'b0;
      13'b0000010000000: n7584_o = 1'b0;
      13'b0000001000000: n7584_o = 1'b0;
      13'b0000000100000: n7584_o = 1'b0;
      13'b0000000010000: n7584_o = 1'b0;
      13'b0000000001000: n7584_o = n6061_o;
      13'b0000000000100: n7584_o = 1'b0;
      13'b0000000000010: n7584_o = 1'b0;
      13'b0000000000001: n7584_o = 1'b0;
      default: n7584_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7586_o = 1'b0;
      13'b0100000000000: n7586_o = n7397_o;
      13'b0010000000000: n7586_o = 1'b0;
      13'b0001000000000: n7586_o = 1'b0;
      13'b0000100000000: n7586_o = 1'b0;
      13'b0000010000000: n7586_o = 1'b0;
      13'b0000001000000: n7586_o = n6459_o;
      13'b0000000100000: n7586_o = 1'b0;
      13'b0000000010000: n7586_o = 1'b0;
      13'b0000000001000: n7586_o = n6062_o;
      13'b0000000000100: n7586_o = n5758_o;
      13'b0000000000010: n7586_o = 1'b0;
      13'b0000000000001: n7586_o = n3083_o;
      default: n7586_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7587_o = n2015_o;
      13'b0100000000000: n7587_o = n2015_o;
      13'b0010000000000: n7587_o = n2015_o;
      13'b0001000000000: n7587_o = n2015_o;
      13'b0000100000000: n7587_o = n2015_o;
      13'b0000010000000: n7587_o = n2015_o;
      13'b0000001000000: n7587_o = n2015_o;
      13'b0000000100000: n7587_o = n2015_o;
      13'b0000000010000: n7587_o = n6125_o;
      13'b0000000001000: n7587_o = n2015_o;
      13'b0000000000100: n7587_o = n5759_o;
      13'b0000000000010: n7587_o = n2015_o;
      13'b0000000000001: n7587_o = n2015_o;
      default: n7587_o = n2015_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7589_o = 1'b0;
      13'b0100000000000: n7589_o = 1'b0;
      13'b0010000000000: n7589_o = 1'b0;
      13'b0001000000000: n7589_o = 1'b0;
      13'b0000100000000: n7589_o = 1'b0;
      13'b0000010000000: n7589_o = 1'b0;
      13'b0000001000000: n7589_o = 1'b0;
      13'b0000000100000: n7589_o = 1'b0;
      13'b0000000010000: n7589_o = n6138_o;
      13'b0000000001000: n7589_o = 1'b0;
      13'b0000000000100: n7589_o = n5761_o;
      13'b0000000000010: n7589_o = 1'b0;
      13'b0000000000001: n7589_o = 1'b0;
      default: n7589_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7591_o = 1'b0;
      13'b0100000000000: n7591_o = 1'b0;
      13'b0010000000000: n7591_o = 1'b0;
      13'b0001000000000: n7591_o = 1'b0;
      13'b0000100000000: n7591_o = 1'b0;
      13'b0000010000000: n7591_o = 1'b0;
      13'b0000001000000: n7591_o = 1'b0;
      13'b0000000100000: n7591_o = 1'b0;
      13'b0000000010000: n7591_o = 1'b0;
      13'b0000000001000: n7591_o = 1'b0;
      13'b0000000000100: n7591_o = n5763_o;
      13'b0000000000010: n7591_o = 1'b0;
      13'b0000000000001: n7591_o = 1'b0;
      default: n7591_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7593_o = 1'b0;
      13'b0100000000000: n7593_o = n7399_o;
      13'b0010000000000: n7593_o = 1'b0;
      13'b0001000000000: n7593_o = 1'b0;
      13'b0000100000000: n7593_o = 1'b0;
      13'b0000010000000: n7593_o = 1'b0;
      13'b0000001000000: n7593_o = 1'b0;
      13'b0000000100000: n7593_o = 1'b0;
      13'b0000000010000: n7593_o = 1'b0;
      13'b0000000001000: n7593_o = 1'b0;
      13'b0000000000100: n7593_o = n5764_o;
      13'b0000000000010: n7593_o = 1'b0;
      13'b0000000000001: n7593_o = 1'b0;
      default: n7593_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7595_o = 1'b0;
      13'b0100000000000: n7595_o = 1'b0;
      13'b0010000000000: n7595_o = n7052_o;
      13'b0001000000000: n7595_o = n6793_o;
      13'b0000100000000: n7595_o = 1'b0;
      13'b0000010000000: n7595_o = n6577_o;
      13'b0000001000000: n7595_o = 1'b0;
      13'b0000000100000: n7595_o = 1'b0;
      13'b0000000010000: n7595_o = 1'b0;
      13'b0000000001000: n7595_o = 1'b0;
      13'b0000000000100: n7595_o = n5765_o;
      13'b0000000000010: n7595_o = n3318_o;
      13'b0000000000001: n7595_o = 1'b0;
      default: n7595_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7597_o = 1'b0;
      13'b0100000000000: n7597_o = n7401_o;
      13'b0010000000000: n7597_o = n7054_o;
      13'b0001000000000: n7597_o = n6795_o;
      13'b0000100000000: n7597_o = 1'b0;
      13'b0000010000000: n7597_o = n6579_o;
      13'b0000001000000: n7597_o = n6460_o;
      13'b0000000100000: n7597_o = 1'b0;
      13'b0000000010000: n7597_o = 1'b0;
      13'b0000000001000: n7597_o = 1'b0;
      13'b0000000000100: n7597_o = n5766_o;
      13'b0000000000010: n7597_o = n3321_o;
      13'b0000000000001: n7597_o = 1'b0;
      default: n7597_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7599_o = 1'b0;
      13'b0100000000000: n7599_o = n7403_o;
      13'b0010000000000: n7599_o = 1'b0;
      13'b0001000000000: n7599_o = 1'b0;
      13'b0000100000000: n7599_o = 1'b0;
      13'b0000010000000: n7599_o = 1'b0;
      13'b0000001000000: n7599_o = 1'b0;
      13'b0000000100000: n7599_o = 1'b0;
      13'b0000000010000: n7599_o = 1'b0;
      13'b0000000001000: n7599_o = 1'b0;
      13'b0000000000100: n7599_o = 1'b0;
      13'b0000000000010: n7599_o = 1'b0;
      13'b0000000000001: n7599_o = 1'b0;
      default: n7599_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7601_o = 1'b0;
      13'b0100000000000: n7601_o = n7405_o;
      13'b0010000000000: n7601_o = 1'b0;
      13'b0001000000000: n7601_o = 1'b0;
      13'b0000100000000: n7601_o = 1'b0;
      13'b0000010000000: n7601_o = 1'b0;
      13'b0000001000000: n7601_o = 1'b0;
      13'b0000000100000: n7601_o = 1'b0;
      13'b0000000010000: n7601_o = 1'b0;
      13'b0000000001000: n7601_o = 1'b0;
      13'b0000000000100: n7601_o = n5768_o;
      13'b0000000000010: n7601_o = 1'b0;
      13'b0000000000001: n7601_o = n3085_o;
      default: n7601_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7603_o = 1'b0;
      13'b0100000000000: n7603_o = 1'b0;
      13'b0010000000000: n7603_o = n7056_o;
      13'b0001000000000: n7603_o = n6797_o;
      13'b0000100000000: n7603_o = 1'b0;
      13'b0000010000000: n7603_o = n6581_o;
      13'b0000001000000: n7603_o = 1'b0;
      13'b0000000100000: n7603_o = 1'b0;
      13'b0000000010000: n7603_o = 1'b0;
      13'b0000000001000: n7603_o = 1'b0;
      13'b0000000000100: n7603_o = n5770_o;
      13'b0000000000010: n7603_o = n3323_o;
      13'b0000000000001: n7603_o = 1'b0;
      default: n7603_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7605_o = 1'b0;
      13'b0100000000000: n7605_o = n7407_o;
      13'b0010000000000: n7605_o = 1'b0;
      13'b0001000000000: n7605_o = 1'b0;
      13'b0000100000000: n7605_o = 1'b0;
      13'b0000010000000: n7605_o = 1'b0;
      13'b0000001000000: n7605_o = 1'b0;
      13'b0000000100000: n7605_o = 1'b0;
      13'b0000000010000: n7605_o = 1'b0;
      13'b0000000001000: n7605_o = 1'b0;
      13'b0000000000100: n7605_o = n5772_o;
      13'b0000000000010: n7605_o = 1'b0;
      13'b0000000000001: n7605_o = 1'b0;
      default: n7605_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7607_o = 1'b0;
      13'b0100000000000: n7607_o = 1'b0;
      13'b0010000000000: n7607_o = n7057_o;
      13'b0001000000000: n7607_o = n6799_o;
      13'b0000100000000: n7607_o = 1'b0;
      13'b0000010000000: n7607_o = n6583_o;
      13'b0000001000000: n7607_o = n6461_o;
      13'b0000000100000: n7607_o = n6156_o;
      13'b0000000010000: n7607_o = 1'b0;
      13'b0000000001000: n7607_o = 1'b0;
      13'b0000000000100: n7607_o = n5773_o;
      13'b0000000000010: n7607_o = n3325_o;
      13'b0000000000001: n7607_o = n3087_o;
      default: n7607_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7608_o = n1900_o;
      13'b0100000000000: n7608_o = n7110_o;
      13'b0010000000000: n7608_o = n1900_o;
      13'b0001000000000: n7608_o = n1900_o;
      13'b0000100000000: n7608_o = n1900_o;
      13'b0000010000000: n7608_o = n1900_o;
      13'b0000001000000: n7608_o = n1900_o;
      13'b0000000100000: n7608_o = n1900_o;
      13'b0000000010000: n7608_o = n1900_o;
      13'b0000000001000: n7608_o = n1900_o;
      13'b0000000000100: n7608_o = n1900_o;
      13'b0000000000010: n7608_o = n1900_o;
      13'b0000000000001: n7608_o = n1900_o;
      default: n7608_o = n1900_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7609_o = n1906_o;
      13'b0100000000000: n7609_o = n1906_o;
      13'b0010000000000: n7609_o = n1906_o;
      13'b0001000000000: n7609_o = n1906_o;
      13'b0000100000000: n7609_o = n1906_o;
      13'b0000010000000: n7609_o = n1906_o;
      13'b0000001000000: n7609_o = n1906_o;
      13'b0000000100000: n7609_o = n1906_o;
      13'b0000000010000: n7609_o = n1906_o;
      13'b0000000001000: n7609_o = n1906_o;
      13'b0000000000100: n7609_o = n5774_o;
      13'b0000000000010: n7609_o = n1906_o;
      13'b0000000000001: n7609_o = n1906_o;
      default: n7609_o = n1906_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7611_o = 1'b0;
      13'b0100000000000: n7611_o = 1'b0;
      13'b0010000000000: n7611_o = 1'b0;
      13'b0001000000000: n7611_o = 1'b0;
      13'b0000100000000: n7611_o = 1'b0;
      13'b0000010000000: n7611_o = 1'b0;
      13'b0000001000000: n7611_o = 1'b0;
      13'b0000000100000: n7611_o = 1'b0;
      13'b0000000010000: n7611_o = 1'b0;
      13'b0000000001000: n7611_o = 1'b0;
      13'b0000000000100: n7611_o = n5776_o;
      13'b0000000000010: n7611_o = 1'b0;
      13'b0000000000001: n7611_o = 1'b0;
      default: n7611_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7612_o = n2154_o;
      13'b0100000000000: n7612_o = n2154_o;
      13'b0010000000000: n7612_o = n2154_o;
      13'b0001000000000: n7612_o = n2154_o;
      13'b0000100000000: n7612_o = n2154_o;
      13'b0000010000000: n7612_o = n2154_o;
      13'b0000001000000: n7612_o = n6462_o;
      13'b0000000100000: n7612_o = n2154_o;
      13'b0000000010000: n7612_o = n2154_o;
      13'b0000000001000: n7612_o = n2154_o;
      13'b0000000000100: n7612_o = n5777_o;
      13'b0000000000010: n7612_o = n2154_o;
      13'b0000000000001: n7612_o = n3088_o;
      default: n7612_o = n2154_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7615_o = n7568_o;
      13'b0100000000000: n7615_o = n7410_o;
      13'b0010000000000: n7615_o = n7058_o;
      13'b0001000000000: n7615_o = n6800_o;
      13'b0000100000000: n7615_o = 1'b0;
      13'b0000010000000: n7615_o = n6586_o;
      13'b0000001000000: n7615_o = n6463_o;
      13'b0000000100000: n7615_o = n6159_o;
      13'b0000000010000: n7615_o = 1'b0;
      13'b0000000001000: n7615_o = n6063_o;
      13'b0000000000100: n7615_o = n5778_o;
      13'b0000000000010: n7615_o = n3328_o;
      13'b0000000000001: n7615_o = n3090_o;
      default: n7615_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7617_o = n7569_o;
      13'b0100000000000: n7617_o = 1'b0;
      13'b0010000000000: n7617_o = 1'b0;
      13'b0001000000000: n7617_o = 1'b0;
      13'b0000100000000: n7617_o = 1'b0;
      13'b0000010000000: n7617_o = 1'b0;
      13'b0000001000000: n7617_o = 1'b0;
      13'b0000000100000: n7617_o = 1'b0;
      13'b0000000010000: n7617_o = 1'b0;
      13'b0000000001000: n7617_o = 1'b0;
      13'b0000000000100: n7617_o = n5780_o;
      13'b0000000000010: n7617_o = 1'b0;
      13'b0000000000001: n7617_o = n3092_o;
      default: n7617_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7620_o = 1'b0;
      13'b0100000000000: n7620_o = 1'b0;
      13'b0010000000000: n7620_o = 1'b0;
      13'b0001000000000: n7620_o = 1'b0;
      13'b0000100000000: n7620_o = 1'b1;
      13'b0000010000000: n7620_o = 1'b0;
      13'b0000001000000: n7620_o = 1'b0;
      13'b0000000100000: n7620_o = 1'b0;
      13'b0000000010000: n7620_o = 1'b0;
      13'b0000000001000: n7620_o = 1'b0;
      13'b0000000000100: n7620_o = 1'b0;
      13'b0000000000010: n7620_o = 1'b0;
      13'b0000000000001: n7620_o = 1'b0;
      default: n7620_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7622_o = n7570_o;
      13'b0100000000000: n7622_o = 1'b0;
      13'b0010000000000: n7622_o = 1'b0;
      13'b0001000000000: n7622_o = 1'b0;
      13'b0000100000000: n7622_o = 1'b0;
      13'b0000010000000: n7622_o = 1'b0;
      13'b0000001000000: n7622_o = 1'b0;
      13'b0000000100000: n7622_o = 1'b0;
      13'b0000000010000: n7622_o = 1'b0;
      13'b0000000001000: n7622_o = 1'b0;
      13'b0000000000100: n7622_o = 1'b0;
      13'b0000000000010: n7622_o = 1'b0;
      13'b0000000000001: n7622_o = 1'b0;
      default: n7622_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7624_o = 1'b0;
      13'b0100000000000: n7624_o = 1'b0;
      13'b0010000000000: n7624_o = 1'b0;
      13'b0001000000000: n7624_o = 1'b0;
      13'b0000100000000: n7624_o = 1'b0;
      13'b0000010000000: n7624_o = 1'b0;
      13'b0000001000000: n7624_o = 1'b0;
      13'b0000000100000: n7624_o = 1'b0;
      13'b0000000010000: n7624_o = 1'b0;
      13'b0000000001000: n7624_o = 1'b0;
      13'b0000000000100: n7624_o = n5782_o;
      13'b0000000000010: n7624_o = 1'b0;
      13'b0000000000001: n7624_o = 1'b0;
      default: n7624_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7626_o = 1'b0;
      13'b0100000000000: n7626_o = 1'b0;
      13'b0010000000000: n7626_o = 1'b0;
      13'b0001000000000: n7626_o = 1'b0;
      13'b0000100000000: n7626_o = 1'b0;
      13'b0000010000000: n7626_o = 1'b0;
      13'b0000001000000: n7626_o = 1'b0;
      13'b0000000100000: n7626_o = 1'b0;
      13'b0000000010000: n7626_o = 1'b0;
      13'b0000000001000: n7626_o = n6065_o;
      13'b0000000000100: n7626_o = n5784_o;
      13'b0000000000010: n7626_o = 1'b0;
      13'b0000000000001: n7626_o = 1'b0;
      default: n7626_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7631_o = 1'b1;
      13'b0100000000000: n7631_o = n7412_o;
      13'b0010000000000: n7631_o = n7059_o;
      13'b0001000000000: n7631_o = n6801_o;
      13'b0000100000000: n7631_o = 1'b1;
      13'b0000010000000: n7631_o = n6589_o;
      13'b0000001000000: n7631_o = n6464_o;
      13'b0000000100000: n7631_o = n6162_o;
      13'b0000000010000: n7631_o = 1'b0;
      13'b0000000001000: n7631_o = n6066_o;
      13'b0000000000100: n7631_o = n5785_o;
      13'b0000000000010: n7631_o = n3331_o;
      13'b0000000000001: n7631_o = n3094_o;
      default: n7631_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7633_o = 1'b0;
      13'b0100000000000: n7633_o = 1'b0;
      13'b0010000000000: n7633_o = 1'b0;
      13'b0001000000000: n7633_o = 1'b0;
      13'b0000100000000: n7633_o = 1'b0;
      13'b0000010000000: n7633_o = 1'b0;
      13'b0000001000000: n7633_o = 1'b0;
      13'b0000000100000: n7633_o = 1'b0;
      13'b0000000010000: n7633_o = 1'b0;
      13'b0000000001000: n7633_o = 1'b0;
      13'b0000000000100: n7633_o = n5787_o;
      13'b0000000000010: n7633_o = 1'b0;
      13'b0000000000001: n7633_o = 1'b0;
      default: n7633_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7635_o = 1'b0;
      13'b0100000000000: n7635_o = n7414_o;
      13'b0010000000000: n7635_o = n7061_o;
      13'b0001000000000: n7635_o = n6802_o;
      13'b0000100000000: n7635_o = 1'b0;
      13'b0000010000000: n7635_o = n6592_o;
      13'b0000001000000: n7635_o = n6466_o;
      13'b0000000100000: n7635_o = 1'b0;
      13'b0000000010000: n7635_o = 1'b0;
      13'b0000000001000: n7635_o = n6067_o;
      13'b0000000000100: n7635_o = n5788_o;
      13'b0000000000010: n7635_o = n3334_o;
      13'b0000000000001: n7635_o = n3096_o;
      default: n7635_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7637_o = 1'b0;
      13'b0100000000000: n7637_o = 1'b0;
      13'b0010000000000: n7637_o = n7063_o;
      13'b0001000000000: n7637_o = n6804_o;
      13'b0000100000000: n7637_o = 1'b0;
      13'b0000010000000: n7637_o = n6594_o;
      13'b0000001000000: n7637_o = n6468_o;
      13'b0000000100000: n7637_o = 1'b0;
      13'b0000000010000: n7637_o = 1'b0;
      13'b0000000001000: n7637_o = 1'b0;
      13'b0000000000100: n7637_o = 1'b0;
      13'b0000000000010: n7637_o = 1'b0;
      13'b0000000000001: n7637_o = 1'b0;
      default: n7637_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7639_o = 1'b0;
      13'b0100000000000: n7639_o = 1'b0;
      13'b0010000000000: n7639_o = n7065_o;
      13'b0001000000000: n7639_o = 1'b0;
      13'b0000100000000: n7639_o = 1'b0;
      13'b0000010000000: n7639_o = n6596_o;
      13'b0000001000000: n7639_o = n6470_o;
      13'b0000000100000: n7639_o = 1'b0;
      13'b0000000010000: n7639_o = 1'b0;
      13'b0000000001000: n7639_o = 1'b0;
      13'b0000000000100: n7639_o = 1'b0;
      13'b0000000000010: n7639_o = 1'b0;
      13'b0000000000001: n7639_o = 1'b0;
      default: n7639_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7641_o = 1'b0;
      13'b0100000000000: n7641_o = 1'b0;
      13'b0010000000000: n7641_o = 1'b0;
      13'b0001000000000: n7641_o = 1'b0;
      13'b0000100000000: n7641_o = 1'b0;
      13'b0000010000000: n7641_o = 1'b0;
      13'b0000001000000: n7641_o = 1'b0;
      13'b0000000100000: n7641_o = 1'b0;
      13'b0000000010000: n7641_o = 1'b0;
      13'b0000000001000: n7641_o = 1'b0;
      13'b0000000000100: n7641_o = 1'b0;
      13'b0000000000010: n7641_o = 1'b0;
      13'b0000000000001: n7641_o = n3098_o;
      default: n7641_o = 1'b0;
    endcase
  assign n7642_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7643_o = n7642_o;
      13'b0100000000000: n7643_o = n7642_o;
      13'b0010000000000: n7643_o = n7642_o;
      13'b0001000000000: n7643_o = n7642_o;
      13'b0000100000000: n7643_o = n7642_o;
      13'b0000010000000: n7643_o = n7642_o;
      13'b0000001000000: n7643_o = n7642_o;
      13'b0000000100000: n7643_o = n7642_o;
      13'b0000000010000: n7643_o = n7642_o;
      13'b0000000001000: n7643_o = n7642_o;
      13'b0000000000100: n7643_o = n5794_o;
      13'b0000000000010: n7643_o = n7642_o;
      13'b0000000000001: n7643_o = n7642_o;
      default: n7643_o = n7642_o;
    endcase
  assign n7644_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7645_o = n7644_o;
      13'b0100000000000: n7645_o = n7644_o;
      13'b0010000000000: n7645_o = n7644_o;
      13'b0001000000000: n7645_o = n7644_o;
      13'b0000100000000: n7645_o = n7644_o;
      13'b0000010000000: n7645_o = n7644_o;
      13'b0000001000000: n7645_o = n7644_o;
      13'b0000000100000: n7645_o = n7644_o;
      13'b0000000010000: n7645_o = n7644_o;
      13'b0000000001000: n7645_o = n7644_o;
      13'b0000000000100: n7645_o = n7644_o;
      13'b0000000000010: n7645_o = n7644_o;
      13'b0000000000001: n7645_o = n3102_o;
      default: n7645_o = n7644_o;
    endcase
  assign n7646_o = n1909_o[20];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7647_o = n7646_o;
      13'b0100000000000: n7647_o = n7646_o;
      13'b0010000000000: n7647_o = n7646_o;
      13'b0001000000000: n7647_o = n7646_o;
      13'b0000100000000: n7647_o = n7646_o;
      13'b0000010000000: n7647_o = n7646_o;
      13'b0000001000000: n7647_o = n7646_o;
      13'b0000000100000: n7647_o = n7646_o;
      13'b0000000010000: n7647_o = n7646_o;
      13'b0000000001000: n7647_o = n7646_o;
      13'b0000000000100: n7647_o = n5796_o;
      13'b0000000000010: n7647_o = n7646_o;
      13'b0000000000001: n7647_o = n7646_o;
      default: n7647_o = n7646_o;
    endcase
  assign n7648_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7649_o = n7648_o;
      13'b0100000000000: n7649_o = n7648_o;
      13'b0010000000000: n7649_o = n7648_o;
      13'b0001000000000: n7649_o = n7648_o;
      13'b0000100000000: n7649_o = n7648_o;
      13'b0000010000000: n7649_o = n7648_o;
      13'b0000001000000: n7649_o = n7648_o;
      13'b0000000100000: n7649_o = n7648_o;
      13'b0000000010000: n7649_o = n7648_o;
      13'b0000000001000: n7649_o = n7648_o;
      13'b0000000000100: n7649_o = n5798_o;
      13'b0000000000010: n7649_o = n7648_o;
      13'b0000000000001: n7649_o = n7648_o;
      default: n7649_o = n7648_o;
    endcase
  assign n7650_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7651_o = n7650_o;
      13'b0100000000000: n7651_o = n7650_o;
      13'b0010000000000: n7651_o = n7650_o;
      13'b0001000000000: n7651_o = n7650_o;
      13'b0000100000000: n7651_o = n7650_o;
      13'b0000010000000: n7651_o = n7650_o;
      13'b0000001000000: n7651_o = n7650_o;
      13'b0000000100000: n7651_o = n7650_o;
      13'b0000000010000: n7651_o = n7650_o;
      13'b0000000001000: n7651_o = n7650_o;
      13'b0000000000100: n7651_o = n7650_o;
      13'b0000000000010: n7651_o = n7650_o;
      13'b0000000000001: n7651_o = n3104_o;
      default: n7651_o = n7650_o;
    endcase
  assign n7652_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7653_o = n7652_o;
      13'b0100000000000: n7653_o = n7416_o;
      13'b0010000000000: n7653_o = n7652_o;
      13'b0001000000000: n7653_o = n7652_o;
      13'b0000100000000: n7653_o = n7652_o;
      13'b0000010000000: n7653_o = n7652_o;
      13'b0000001000000: n7653_o = n7652_o;
      13'b0000000100000: n7653_o = n7652_o;
      13'b0000000010000: n7653_o = n7652_o;
      13'b0000000001000: n7653_o = n7652_o;
      13'b0000000000100: n7653_o = n7652_o;
      13'b0000000000010: n7653_o = n7652_o;
      13'b0000000000001: n7653_o = n7652_o;
      default: n7653_o = n7652_o;
    endcase
  assign n7654_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7655_o = n7654_o;
      13'b0100000000000: n7655_o = n7654_o;
      13'b0010000000000: n7655_o = n7067_o;
      13'b0001000000000: n7655_o = n7654_o;
      13'b0000100000000: n7655_o = n7654_o;
      13'b0000010000000: n7655_o = n7654_o;
      13'b0000001000000: n7655_o = n7654_o;
      13'b0000000100000: n7655_o = n7654_o;
      13'b0000000010000: n7655_o = n7654_o;
      13'b0000000001000: n7655_o = n7654_o;
      13'b0000000000100: n7655_o = n5800_o;
      13'b0000000000010: n7655_o = n7654_o;
      13'b0000000000001: n7655_o = n7654_o;
      default: n7655_o = n7654_o;
    endcase
  assign n7656_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7657_o = n7656_o;
      13'b0100000000000: n7657_o = n7656_o;
      13'b0010000000000: n7657_o = n7656_o;
      13'b0001000000000: n7657_o = n7656_o;
      13'b0000100000000: n7657_o = n7656_o;
      13'b0000010000000: n7657_o = n7656_o;
      13'b0000001000000: n7657_o = n7656_o;
      13'b0000000100000: n7657_o = n7656_o;
      13'b0000000010000: n7657_o = n7656_o;
      13'b0000000001000: n7657_o = n7656_o;
      13'b0000000000100: n7657_o = n5802_o;
      13'b0000000000010: n7657_o = n7656_o;
      13'b0000000000001: n7657_o = n7656_o;
      default: n7657_o = n7656_o;
    endcase
  assign n7658_o = n1909_o[37];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7659_o = n7658_o;
      13'b0100000000000: n7659_o = n7658_o;
      13'b0010000000000: n7659_o = n7658_o;
      13'b0001000000000: n7659_o = n7658_o;
      13'b0000100000000: n7659_o = n7658_o;
      13'b0000010000000: n7659_o = n7658_o;
      13'b0000001000000: n7659_o = n7658_o;
      13'b0000000100000: n7659_o = n7658_o;
      13'b0000000010000: n7659_o = n7658_o;
      13'b0000000001000: n7659_o = n7658_o;
      13'b0000000000100: n7659_o = n7658_o;
      13'b0000000000010: n7659_o = n7658_o;
      13'b0000000000001: n7659_o = n3106_o;
      default: n7659_o = n7658_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7660_o = n2007_o;
      13'b0100000000000: n7660_o = n2007_o;
      13'b0010000000000: n7660_o = n2007_o;
      13'b0001000000000: n7660_o = n6805_o;
      13'b0000100000000: n7660_o = n2007_o;
      13'b0000010000000: n7660_o = n2007_o;
      13'b0000001000000: n7660_o = n2007_o;
      13'b0000000100000: n7660_o = n2007_o;
      13'b0000000010000: n7660_o = n2007_o;
      13'b0000000001000: n7660_o = n2007_o;
      13'b0000000000100: n7660_o = n2007_o;
      13'b0000000000010: n7660_o = n2007_o;
      13'b0000000000001: n7660_o = n2007_o;
      default: n7660_o = n2007_o;
    endcase
  assign n7661_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7662_o = n7661_o;
      13'b0100000000000: n7662_o = n7661_o;
      13'b0010000000000: n7662_o = n7661_o;
      13'b0001000000000: n7662_o = n7661_o;
      13'b0000100000000: n7662_o = n7661_o;
      13'b0000010000000: n7662_o = n7661_o;
      13'b0000001000000: n7662_o = n7661_o;
      13'b0000000100000: n7662_o = n7661_o;
      13'b0000000010000: n7662_o = n7661_o;
      13'b0000000001000: n7662_o = n7661_o;
      13'b0000000000100: n7662_o = n7661_o;
      13'b0000000000010: n7662_o = n7661_o;
      13'b0000000000001: n7662_o = n3108_o;
      default: n7662_o = n7661_o;
    endcase
  assign n7663_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7664_o = n7663_o;
      13'b0100000000000: n7664_o = n7663_o;
      13'b0010000000000: n7664_o = n7663_o;
      13'b0001000000000: n7664_o = n7663_o;
      13'b0000100000000: n7664_o = n7663_o;
      13'b0000010000000: n7664_o = n7663_o;
      13'b0000001000000: n7664_o = n7663_o;
      13'b0000000100000: n7664_o = n7663_o;
      13'b0000000010000: n7664_o = n7663_o;
      13'b0000000001000: n7664_o = n7663_o;
      13'b0000000000100: n7664_o = n5804_o;
      13'b0000000000010: n7664_o = n3308_o;
      13'b0000000000001: n7664_o = n7663_o;
      default: n7664_o = n7663_o;
    endcase
  assign n7665_o = n3110_o[0];
  assign n7666_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7667_o = n7666_o;
      13'b0100000000000: n7667_o = n7418_o;
      13'b0010000000000: n7667_o = n7666_o;
      13'b0001000000000: n7667_o = n7666_o;
      13'b0000100000000: n7667_o = n7666_o;
      13'b0000010000000: n7667_o = n7666_o;
      13'b0000001000000: n7667_o = n7666_o;
      13'b0000000100000: n7667_o = n7666_o;
      13'b0000000010000: n7667_o = n7666_o;
      13'b0000000001000: n7667_o = n7666_o;
      13'b0000000000100: n7667_o = n5806_o;
      13'b0000000000010: n7667_o = n7666_o;
      13'b0000000000001: n7667_o = n7665_o;
      default: n7667_o = n7666_o;
    endcase
  assign n7668_o = n3110_o[1];
  assign n7669_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7670_o = n7669_o;
      13'b0100000000000: n7670_o = n7669_o;
      13'b0010000000000: n7670_o = n7669_o;
      13'b0001000000000: n7670_o = n7669_o;
      13'b0000100000000: n7670_o = n7669_o;
      13'b0000010000000: n7670_o = n7669_o;
      13'b0000001000000: n7670_o = n7669_o;
      13'b0000000100000: n7670_o = n7669_o;
      13'b0000000010000: n7670_o = n7669_o;
      13'b0000000001000: n7670_o = n7669_o;
      13'b0000000000100: n7670_o = n5808_o;
      13'b0000000000010: n7670_o = n7669_o;
      13'b0000000000001: n7670_o = n7668_o;
      default: n7670_o = n7669_o;
    endcase
  assign n7671_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7672_o = n7671_o;
      13'b0100000000000: n7672_o = n7671_o;
      13'b0010000000000: n7672_o = n7671_o;
      13'b0001000000000: n7672_o = n7671_o;
      13'b0000100000000: n7672_o = n7671_o;
      13'b0000010000000: n7672_o = n7671_o;
      13'b0000001000000: n7672_o = n6472_o;
      13'b0000000100000: n7672_o = n7671_o;
      13'b0000000010000: n7672_o = n7671_o;
      13'b0000000001000: n7672_o = n7671_o;
      13'b0000000000100: n7672_o = n5810_o;
      13'b0000000000010: n7672_o = n7671_o;
      13'b0000000000001: n7672_o = n7671_o;
      default: n7672_o = n7671_o;
    endcase
  assign n7673_o = n3309_o[0];
  assign n7674_o = n5814_o[0];
  assign n7675_o = n2162_o[0];
  assign n7676_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n7677_o = n2037_o ? n7675_o : n7676_o;
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7678_o = n7677_o;
      13'b0100000000000: n7678_o = n7677_o;
      13'b0010000000000: n7678_o = n7677_o;
      13'b0001000000000: n7678_o = n6809_o;
      13'b0000100000000: n7678_o = n7677_o;
      13'b0000010000000: n7678_o = n7677_o;
      13'b0000001000000: n7678_o = n7677_o;
      13'b0000000100000: n7678_o = n7677_o;
      13'b0000000010000: n7678_o = n7677_o;
      13'b0000000001000: n7678_o = n7677_o;
      13'b0000000000100: n7678_o = n7674_o;
      13'b0000000000010: n7678_o = n7673_o;
      13'b0000000000001: n7678_o = n7677_o;
      default: n7678_o = n7677_o;
    endcase
  assign n7679_o = n3309_o[1];
  assign n7680_o = n5814_o[1];
  assign n7681_o = n2162_o[1];
  assign n7682_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n7683_o = n2037_o ? n7681_o : n7682_o;
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7684_o = n7683_o;
      13'b0100000000000: n7684_o = n7683_o;
      13'b0010000000000: n7684_o = n7683_o;
      13'b0001000000000: n7684_o = n7683_o;
      13'b0000100000000: n7684_o = n7683_o;
      13'b0000010000000: n7684_o = n7683_o;
      13'b0000001000000: n7684_o = n7683_o;
      13'b0000000100000: n7684_o = n7683_o;
      13'b0000000010000: n7684_o = n6142_o;
      13'b0000000001000: n7684_o = n7683_o;
      13'b0000000000100: n7684_o = n7680_o;
      13'b0000000000010: n7684_o = n7679_o;
      13'b0000000000001: n7684_o = n7683_o;
      default: n7684_o = n7683_o;
    endcase
  assign n7685_o = n5814_o[2];
  assign n7686_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7687_o = n7686_o;
      13'b0100000000000: n7687_o = n7686_o;
      13'b0010000000000: n7687_o = n7686_o;
      13'b0001000000000: n7687_o = n7686_o;
      13'b0000100000000: n7687_o = n7686_o;
      13'b0000010000000: n7687_o = n7686_o;
      13'b0000001000000: n7687_o = n7686_o;
      13'b0000000100000: n7687_o = n7686_o;
      13'b0000000010000: n7687_o = n7686_o;
      13'b0000000001000: n7687_o = n7686_o;
      13'b0000000000100: n7687_o = n7685_o;
      13'b0000000000010: n7687_o = n7686_o;
      13'b0000000000001: n7687_o = n7686_o;
      default: n7687_o = n7686_o;
    endcase
  assign n7688_o = n3341_o[0];
  assign n7689_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7690_o = n7689_o;
      13'b0100000000000: n7690_o = n7689_o;
      13'b0010000000000: n7690_o = n7689_o;
      13'b0001000000000: n7690_o = n7689_o;
      13'b0000100000000: n7690_o = n7689_o;
      13'b0000010000000: n7690_o = n6572_o;
      13'b0000001000000: n7690_o = n6474_o;
      13'b0000000100000: n7690_o = n7689_o;
      13'b0000000010000: n7690_o = n7689_o;
      13'b0000000001000: n7690_o = n6069_o;
      13'b0000000000100: n7690_o = n5816_o;
      13'b0000000000010: n7690_o = n7688_o;
      13'b0000000000001: n7690_o = n3112_o;
      default: n7690_o = n7689_o;
    endcase
  assign n7691_o = n3341_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7692_o = n2168_o;
      13'b0100000000000: n7692_o = n2168_o;
      13'b0010000000000: n7692_o = n2168_o;
      13'b0001000000000: n7692_o = n6810_o;
      13'b0000100000000: n7692_o = n2168_o;
      13'b0000010000000: n7692_o = n2168_o;
      13'b0000001000000: n7692_o = n2168_o;
      13'b0000000100000: n7692_o = n2168_o;
      13'b0000000010000: n7692_o = n2168_o;
      13'b0000000001000: n7692_o = n2168_o;
      13'b0000000000100: n7692_o = n2168_o;
      13'b0000000000010: n7692_o = n7691_o;
      13'b0000000000001: n7692_o = n3114_o;
      default: n7692_o = n2168_o;
    endcase
  assign n7693_o = n5819_o[1:0];
  assign n7694_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7695_o = n7694_o;
      13'b0100000000000: n7695_o = n7694_o;
      13'b0010000000000: n7695_o = n7694_o;
      13'b0001000000000: n7695_o = n7694_o;
      13'b0000100000000: n7695_o = n7694_o;
      13'b0000010000000: n7695_o = n7694_o;
      13'b0000001000000: n7695_o = n7694_o;
      13'b0000000100000: n7695_o = n7694_o;
      13'b0000000010000: n7695_o = n7694_o;
      13'b0000000001000: n7695_o = n7694_o;
      13'b0000000000100: n7695_o = n7693_o;
      13'b0000000000010: n7695_o = n7694_o;
      13'b0000000000001: n7695_o = n3116_o;
      default: n7695_o = n7694_o;
    endcase
  assign n7696_o = n5819_o[2];
  assign n7697_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7698_o = n7697_o;
      13'b0100000000000: n7698_o = n7697_o;
      13'b0010000000000: n7698_o = n7697_o;
      13'b0001000000000: n7698_o = n7697_o;
      13'b0000100000000: n7698_o = n7697_o;
      13'b0000010000000: n7698_o = n7697_o;
      13'b0000001000000: n7698_o = n7697_o;
      13'b0000000100000: n7698_o = n7697_o;
      13'b0000000010000: n7698_o = n7697_o;
      13'b0000000001000: n7698_o = n5876_o;
      13'b0000000000100: n7698_o = n7696_o;
      13'b0000000000010: n7698_o = n7697_o;
      13'b0000000000001: n7698_o = n7697_o;
      default: n7698_o = n7697_o;
    endcase
  assign n7699_o = n5819_o[3];
  assign n7700_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7701_o = n7700_o;
      13'b0100000000000: n7701_o = n7700_o;
      13'b0010000000000: n7701_o = n7700_o;
      13'b0001000000000: n7701_o = n7700_o;
      13'b0000100000000: n7701_o = n7700_o;
      13'b0000010000000: n7701_o = n7700_o;
      13'b0000001000000: n7701_o = n7700_o;
      13'b0000000100000: n7701_o = n7700_o;
      13'b0000000010000: n7701_o = n7700_o;
      13'b0000000001000: n7701_o = n7700_o;
      13'b0000000000100: n7701_o = n7699_o;
      13'b0000000000010: n7701_o = n7700_o;
      13'b0000000000001: n7701_o = n7700_o;
      default: n7701_o = n7700_o;
    endcase
  assign n7702_o = n3118_o[0];
  assign n7703_o = n5819_o[4];
  assign n7704_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7705_o = n7704_o;
      13'b0100000000000: n7705_o = n7420_o;
      13'b0010000000000: n7705_o = n7704_o;
      13'b0001000000000: n7705_o = n7704_o;
      13'b0000100000000: n7705_o = n7704_o;
      13'b0000010000000: n7705_o = n7704_o;
      13'b0000001000000: n7705_o = n7704_o;
      13'b0000000100000: n7705_o = n7704_o;
      13'b0000000010000: n7705_o = n7704_o;
      13'b0000000001000: n7705_o = n7704_o;
      13'b0000000000100: n7705_o = n7703_o;
      13'b0000000000010: n7705_o = n7704_o;
      13'b0000000000001: n7705_o = n7702_o;
      default: n7705_o = n7704_o;
    endcase
  assign n7706_o = n3118_o[1];
  assign n7707_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7708_o = n7707_o;
      13'b0100000000000: n7708_o = n7707_o;
      13'b0010000000000: n7708_o = n7707_o;
      13'b0001000000000: n7708_o = n6811_o;
      13'b0000100000000: n7708_o = n7707_o;
      13'b0000010000000: n7708_o = n6526_o;
      13'b0000001000000: n7708_o = n6476_o;
      13'b0000000100000: n7708_o = n7707_o;
      13'b0000000010000: n7708_o = n7707_o;
      13'b0000000001000: n7708_o = n6073_o;
      13'b0000000000100: n7708_o = n5821_o;
      13'b0000000000010: n7708_o = n7707_o;
      13'b0000000000001: n7708_o = n7706_o;
      default: n7708_o = n7707_o;
    endcase
  assign n7709_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7710_o = n7709_o;
      13'b0100000000000: n7710_o = n7709_o;
      13'b0010000000000: n7710_o = n7709_o;
      13'b0001000000000: n7710_o = n7709_o;
      13'b0000100000000: n7710_o = n7709_o;
      13'b0000010000000: n7710_o = n7709_o;
      13'b0000001000000: n7710_o = n7709_o;
      13'b0000000100000: n7710_o = n7709_o;
      13'b0000000010000: n7710_o = n7709_o;
      13'b0000000001000: n7710_o = n7709_o;
      13'b0000000000100: n7710_o = n5824_o;
      13'b0000000000010: n7710_o = n7709_o;
      13'b0000000000001: n7710_o = n7709_o;
      default: n7710_o = n7709_o;
    endcase
  assign n7711_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7712_o = n7711_o;
      13'b0100000000000: n7712_o = n7711_o;
      13'b0010000000000: n7712_o = n7069_o;
      13'b0001000000000: n7712_o = n7711_o;
      13'b0000100000000: n7712_o = n7711_o;
      13'b0000010000000: n7712_o = n7711_o;
      13'b0000001000000: n7712_o = n7711_o;
      13'b0000000100000: n7712_o = n7711_o;
      13'b0000000010000: n7712_o = n7711_o;
      13'b0000000001000: n7712_o = n7711_o;
      13'b0000000000100: n7712_o = n7711_o;
      13'b0000000000010: n7712_o = n7711_o;
      13'b0000000000001: n7712_o = n7711_o;
      default: n7712_o = n7711_o;
    endcase
  assign n7713_o = n1909_o[67];
  assign n7714_o = {n7713_o, n2019_o, n2178_o};
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7715_o = n7714_o;
      13'b0100000000000: n7715_o = n7714_o;
      13'b0010000000000: n7715_o = n7714_o;
      13'b0001000000000: n7715_o = n7714_o;
      13'b0000100000000: n7715_o = n7714_o;
      13'b0000010000000: n7715_o = n7714_o;
      13'b0000001000000: n7715_o = n7714_o;
      13'b0000000100000: n7715_o = n7714_o;
      13'b0000000010000: n7715_o = n7714_o;
      13'b0000000001000: n7715_o = n7714_o;
      13'b0000000000100: n7715_o = n5827_o;
      13'b0000000000010: n7715_o = n7714_o;
      13'b0000000000001: n7715_o = n7714_o;
      default: n7715_o = n7714_o;
    endcase
  assign n7716_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7717_o = n7716_o;
      13'b0100000000000: n7717_o = n7716_o;
      13'b0010000000000: n7717_o = n7716_o;
      13'b0001000000000: n7717_o = n7716_o;
      13'b0000100000000: n7717_o = n7716_o;
      13'b0000010000000: n7717_o = n7716_o;
      13'b0000001000000: n7717_o = n7716_o;
      13'b0000000100000: n7717_o = n7716_o;
      13'b0000000010000: n7717_o = n7716_o;
      13'b0000000001000: n7717_o = n7716_o;
      13'b0000000000100: n7717_o = n5829_o;
      13'b0000000000010: n7717_o = n7716_o;
      13'b0000000000001: n7717_o = n7716_o;
      default: n7717_o = n7716_o;
    endcase
  assign n7718_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7719_o = n7718_o;
      13'b0100000000000: n7719_o = n7422_o;
      13'b0010000000000: n7719_o = n7718_o;
      13'b0001000000000: n7719_o = n7718_o;
      13'b0000100000000: n7719_o = n7718_o;
      13'b0000010000000: n7719_o = n7718_o;
      13'b0000001000000: n7719_o = n7718_o;
      13'b0000000100000: n7719_o = n7718_o;
      13'b0000000010000: n7719_o = n7718_o;
      13'b0000000001000: n7719_o = n7718_o;
      13'b0000000000100: n7719_o = n5831_o;
      13'b0000000000010: n7719_o = n7718_o;
      13'b0000000000001: n7719_o = n3120_o;
      default: n7719_o = n7718_o;
    endcase
  assign n7720_o = n5834_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7721_o = n2171_o;
      13'b0100000000000: n7721_o = n2171_o;
      13'b0010000000000: n7721_o = n2171_o;
      13'b0001000000000: n7721_o = n2171_o;
      13'b0000100000000: n7721_o = n2171_o;
      13'b0000010000000: n7721_o = n2171_o;
      13'b0000001000000: n7721_o = n2171_o;
      13'b0000000100000: n7721_o = n2171_o;
      13'b0000000010000: n7721_o = n6143_o;
      13'b0000000001000: n7721_o = n6074_o;
      13'b0000000000100: n7721_o = n7720_o;
      13'b0000000000010: n7721_o = n3311_o;
      13'b0000000000001: n7721_o = n3121_o;
      default: n7721_o = n2171_o;
    endcase
  assign n7722_o = n5834_o[1];
  assign n7723_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7724_o = n7723_o;
      13'b0100000000000: n7724_o = n7723_o;
      13'b0010000000000: n7724_o = n7723_o;
      13'b0001000000000: n7724_o = n7723_o;
      13'b0000100000000: n7724_o = n7723_o;
      13'b0000010000000: n7724_o = n7723_o;
      13'b0000001000000: n7724_o = n7723_o;
      13'b0000000100000: n7724_o = n7723_o;
      13'b0000000010000: n7724_o = n7723_o;
      13'b0000000001000: n7724_o = n7723_o;
      13'b0000000000100: n7724_o = n7722_o;
      13'b0000000000010: n7724_o = n7723_o;
      13'b0000000000001: n7724_o = n7723_o;
      default: n7724_o = n7723_o;
    endcase
  assign n7725_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7726_o = n7725_o;
      13'b0100000000000: n7726_o = n7725_o;
      13'b0010000000000: n7726_o = n7725_o;
      13'b0001000000000: n7726_o = n7725_o;
      13'b0000100000000: n7726_o = n7725_o;
      13'b0000010000000: n7726_o = n7725_o;
      13'b0000001000000: n7726_o = n6478_o;
      13'b0000000100000: n7726_o = n7725_o;
      13'b0000000010000: n7726_o = n7725_o;
      13'b0000000001000: n7726_o = n7725_o;
      13'b0000000000100: n7726_o = n7725_o;
      13'b0000000000010: n7726_o = n7725_o;
      13'b0000000000001: n7726_o = n7725_o;
      default: n7726_o = n7725_o;
    endcase
  assign n7727_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7728_o = n7727_o;
      13'b0100000000000: n7728_o = n7727_o;
      13'b0010000000000: n7728_o = n7727_o;
      13'b0001000000000: n7728_o = n7727_o;
      13'b0000100000000: n7728_o = n7727_o;
      13'b0000010000000: n7728_o = n7727_o;
      13'b0000001000000: n7728_o = n7727_o;
      13'b0000000100000: n7728_o = n7727_o;
      13'b0000000010000: n7728_o = n7727_o;
      13'b0000000001000: n7728_o = n7727_o;
      13'b0000000000100: n7728_o = n7727_o;
      13'b0000000000010: n7728_o = n7727_o;
      13'b0000000000001: n7728_o = n3123_o;
      default: n7728_o = n7727_o;
    endcase
  assign n7729_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7730_o = n7729_o;
      13'b0100000000000: n7730_o = n7729_o;
      13'b0010000000000: n7730_o = n7729_o;
      13'b0001000000000: n7730_o = n7729_o;
      13'b0000100000000: n7730_o = n7729_o;
      13'b0000010000000: n7730_o = n7729_o;
      13'b0000001000000: n7730_o = n7729_o;
      13'b0000000100000: n7730_o = n7729_o;
      13'b0000000010000: n7730_o = n7729_o;
      13'b0000000001000: n7730_o = n7729_o;
      13'b0000000000100: n7730_o = n7729_o;
      13'b0000000000010: n7730_o = n7729_o;
      13'b0000000000001: n7730_o = n3125_o;
      default: n7730_o = n7729_o;
    endcase
  assign n7731_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7732_o = n7731_o;
      13'b0100000000000: n7732_o = n7731_o;
      13'b0010000000000: n7732_o = n7071_o;
      13'b0001000000000: n7732_o = n7731_o;
      13'b0000100000000: n7732_o = n7731_o;
      13'b0000010000000: n7732_o = n7731_o;
      13'b0000001000000: n7732_o = n7731_o;
      13'b0000000100000: n7732_o = n7731_o;
      13'b0000000010000: n7732_o = n7731_o;
      13'b0000000001000: n7732_o = n7731_o;
      13'b0000000000100: n7732_o = n7731_o;
      13'b0000000000010: n7732_o = n7731_o;
      13'b0000000000001: n7732_o = n7731_o;
      default: n7732_o = n7731_o;
    endcase
  assign n7733_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7734_o = n7733_o;
      13'b0100000000000: n7734_o = n7733_o;
      13'b0010000000000: n7734_o = n7733_o;
      13'b0001000000000: n7734_o = n7733_o;
      13'b0000100000000: n7734_o = n7733_o;
      13'b0000010000000: n7734_o = n7733_o;
      13'b0000001000000: n7734_o = n7733_o;
      13'b0000000100000: n7734_o = n7733_o;
      13'b0000000010000: n7734_o = n7733_o;
      13'b0000000001000: n7734_o = n7733_o;
      13'b0000000000100: n7734_o = n7733_o;
      13'b0000000000010: n7734_o = n7733_o;
      13'b0000000000001: n7734_o = n3127_o;
      default: n7734_o = n7733_o;
    endcase
  assign n7735_o = n6165_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7737_o = 1'b0;
      13'b0100000000000: n7737_o = 1'b0;
      13'b0010000000000: n7737_o = 1'b0;
      13'b0001000000000: n7737_o = 1'b0;
      13'b0000100000000: n7737_o = 1'b0;
      13'b0000010000000: n7737_o = 1'b0;
      13'b0000001000000: n7737_o = 1'b0;
      13'b0000000100000: n7737_o = n7735_o;
      13'b0000000010000: n7737_o = 1'b0;
      13'b0000000001000: n7737_o = 1'b0;
      13'b0000000000100: n7737_o = n5838_o;
      13'b0000000000010: n7737_o = n3344_o;
      13'b0000000000001: n7737_o = n3129_o;
      default: n7737_o = 1'b0;
    endcase
  assign n7738_o = n6165_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7740_o = 1'b0;
      13'b0100000000000: n7740_o = 1'b0;
      13'b0010000000000: n7740_o = 1'b0;
      13'b0001000000000: n7740_o = 1'b0;
      13'b0000100000000: n7740_o = 1'b0;
      13'b0000010000000: n7740_o = 1'b0;
      13'b0000001000000: n7740_o = 1'b0;
      13'b0000000100000: n7740_o = n7738_o;
      13'b0000000010000: n7740_o = 1'b0;
      13'b0000000001000: n7740_o = 1'b0;
      13'b0000000000100: n7740_o = 1'b0;
      13'b0000000000010: n7740_o = 1'b0;
      13'b0000000000001: n7740_o = 1'b0;
      default: n7740_o = 1'b0;
    endcase
  assign n7741_o = n5840_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7743_o = 1'b0;
      13'b0100000000000: n7743_o = 1'b0;
      13'b0010000000000: n7743_o = 1'b0;
      13'b0001000000000: n7743_o = 1'b0;
      13'b0000100000000: n7743_o = 1'b0;
      13'b0000010000000: n7743_o = 1'b0;
      13'b0000001000000: n7743_o = 1'b0;
      13'b0000000100000: n7743_o = 1'b0;
      13'b0000000010000: n7743_o = 1'b0;
      13'b0000000001000: n7743_o = 1'b0;
      13'b0000000000100: n7743_o = n7741_o;
      13'b0000000000010: n7743_o = 1'b0;
      13'b0000000000001: n7743_o = 1'b0;
      default: n7743_o = 1'b0;
    endcase
  assign n7744_o = n5840_o[1];
  assign n7745_o = n6076_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7747_o = 1'b0;
      13'b0100000000000: n7747_o = 1'b0;
      13'b0010000000000: n7747_o = n7073_o;
      13'b0001000000000: n7747_o = 1'b0;
      13'b0000100000000: n7747_o = 1'b0;
      13'b0000010000000: n7747_o = n6602_o;
      13'b0000001000000: n7747_o = n6480_o;
      13'b0000000100000: n7747_o = 1'b0;
      13'b0000000010000: n7747_o = 1'b0;
      13'b0000000001000: n7747_o = n7745_o;
      13'b0000000000100: n7747_o = n7744_o;
      13'b0000000000010: n7747_o = 1'b0;
      13'b0000000000001: n7747_o = n3131_o;
      default: n7747_o = 1'b0;
    endcase
  assign n7748_o = n6076_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7750_o = 1'b0;
      13'b0100000000000: n7750_o = 1'b0;
      13'b0010000000000: n7750_o = 1'b0;
      13'b0001000000000: n7750_o = 1'b0;
      13'b0000100000000: n7750_o = 1'b0;
      13'b0000010000000: n7750_o = 1'b0;
      13'b0000001000000: n7750_o = 1'b0;
      13'b0000000100000: n7750_o = 1'b0;
      13'b0000000010000: n7750_o = 1'b0;
      13'b0000000001000: n7750_o = n7748_o;
      13'b0000000000100: n7750_o = 1'b0;
      13'b0000000000010: n7750_o = 1'b0;
      13'b0000000000001: n7750_o = 1'b0;
      default: n7750_o = 1'b0;
    endcase
  assign n7751_o = n3133_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7753_o = 1'b0;
      13'b0100000000000: n7753_o = 1'b0;
      13'b0010000000000: n7753_o = 1'b0;
      13'b0001000000000: n7753_o = 1'b0;
      13'b0000100000000: n7753_o = 1'b0;
      13'b0000010000000: n7753_o = 1'b0;
      13'b0000001000000: n7753_o = n6482_o;
      13'b0000000100000: n7753_o = 1'b0;
      13'b0000000010000: n7753_o = 1'b0;
      13'b0000000001000: n7753_o = 1'b0;
      13'b0000000000100: n7753_o = 1'b0;
      13'b0000000000010: n7753_o = 1'b0;
      13'b0000000000001: n7753_o = n7751_o;
      default: n7753_o = 1'b0;
    endcase
  assign n7754_o = n3133_o[1];
  assign n7755_o = n5842_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7757_o = 1'b0;
      13'b0100000000000: n7757_o = 1'b0;
      13'b0010000000000: n7757_o = n7075_o;
      13'b0001000000000: n7757_o = 1'b0;
      13'b0000100000000: n7757_o = 1'b0;
      13'b0000010000000: n7757_o = 1'b0;
      13'b0000001000000: n7757_o = 1'b0;
      13'b0000000100000: n7757_o = 1'b0;
      13'b0000000010000: n7757_o = 1'b0;
      13'b0000000001000: n7757_o = 1'b0;
      13'b0000000000100: n7757_o = n7755_o;
      13'b0000000000010: n7757_o = 1'b0;
      13'b0000000000001: n7757_o = n7754_o;
      default: n7757_o = 1'b0;
    endcase
  assign n7758_o = n3133_o[2];
  assign n7759_o = n5842_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7761_o = 1'b0;
      13'b0100000000000: n7761_o = 1'b0;
      13'b0010000000000: n7761_o = 1'b0;
      13'b0001000000000: n7761_o = n6815_o;
      13'b0000100000000: n7761_o = 1'b0;
      13'b0000010000000: n7761_o = 1'b0;
      13'b0000001000000: n7761_o = 1'b0;
      13'b0000000100000: n7761_o = 1'b0;
      13'b0000000010000: n7761_o = 1'b0;
      13'b0000000001000: n7761_o = 1'b0;
      13'b0000000000100: n7761_o = n7759_o;
      13'b0000000000010: n7761_o = 1'b0;
      13'b0000000000001: n7761_o = n7758_o;
      default: n7761_o = 1'b0;
    endcase
  assign n7762_o = n3133_o[3];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7764_o = 1'b0;
      13'b0100000000000: n7764_o = 1'b0;
      13'b0010000000000: n7764_o = 1'b0;
      13'b0001000000000: n7764_o = n6817_o;
      13'b0000100000000: n7764_o = 1'b0;
      13'b0000010000000: n7764_o = 1'b0;
      13'b0000001000000: n7764_o = 1'b0;
      13'b0000000100000: n7764_o = 1'b0;
      13'b0000000010000: n7764_o = 1'b0;
      13'b0000000001000: n7764_o = 1'b0;
      13'b0000000000100: n7764_o = 1'b0;
      13'b0000000000010: n7764_o = 1'b0;
      13'b0000000000001: n7764_o = n7762_o;
      default: n7764_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7766_o = 1'b0;
      13'b0100000000000: n7766_o = 1'b0;
      13'b0010000000000: n7766_o = 1'b0;
      13'b0001000000000: n7766_o = n6819_o;
      13'b0000100000000: n7766_o = 1'b0;
      13'b0000010000000: n7766_o = 1'b0;
      13'b0000001000000: n7766_o = 1'b0;
      13'b0000000100000: n7766_o = 1'b0;
      13'b0000000010000: n7766_o = 1'b0;
      13'b0000000001000: n7766_o = 1'b0;
      13'b0000000000100: n7766_o = 1'b0;
      13'b0000000000010: n7766_o = 1'b0;
      13'b0000000000001: n7766_o = 1'b0;
      default: n7766_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7768_o = 1'b0;
      13'b0100000000000: n7768_o = 1'b0;
      13'b0010000000000: n7768_o = 1'b0;
      13'b0001000000000: n7768_o = 1'b0;
      13'b0000100000000: n7768_o = 1'b0;
      13'b0000010000000: n7768_o = 1'b0;
      13'b0000001000000: n7768_o = 1'b0;
      13'b0000000100000: n7768_o = 1'b0;
      13'b0000000010000: n7768_o = 1'b0;
      13'b0000000001000: n7768_o = 1'b0;
      13'b0000000000100: n7768_o = n5843_o;
      13'b0000000000010: n7768_o = 1'b0;
      13'b0000000000001: n7768_o = 1'b0;
      default: n7768_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7770_o = 1'b0;
      13'b0100000000000: n7770_o = 1'b0;
      13'b0010000000000: n7770_o = n7077_o;
      13'b0001000000000: n7770_o = 1'b0;
      13'b0000100000000: n7770_o = 1'b0;
      13'b0000010000000: n7770_o = 1'b0;
      13'b0000001000000: n7770_o = 1'b0;
      13'b0000000100000: n7770_o = 1'b0;
      13'b0000000010000: n7770_o = 1'b0;
      13'b0000000001000: n7770_o = 1'b0;
      13'b0000000000100: n7770_o = 1'b0;
      13'b0000000000010: n7770_o = 1'b0;
      13'b0000000000001: n7770_o = 1'b0;
      default: n7770_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7772_o = 1'b0;
      13'b0100000000000: n7772_o = 1'b0;
      13'b0010000000000: n7772_o = 1'b0;
      13'b0001000000000: n7772_o = 1'b0;
      13'b0000100000000: n7772_o = 1'b0;
      13'b0000010000000: n7772_o = 1'b0;
      13'b0000001000000: n7772_o = n6484_o;
      13'b0000000100000: n7772_o = 1'b0;
      13'b0000000010000: n7772_o = 1'b0;
      13'b0000000001000: n7772_o = 1'b0;
      13'b0000000000100: n7772_o = n5845_o;
      13'b0000000000010: n7772_o = 1'b0;
      13'b0000000000001: n7772_o = 1'b0;
      default: n7772_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7774_o = 1'b0;
      13'b0100000000000: n7774_o = 1'b0;
      13'b0010000000000: n7774_o = 1'b0;
      13'b0001000000000: n7774_o = 1'b0;
      13'b0000100000000: n7774_o = 1'b0;
      13'b0000010000000: n7774_o = 1'b0;
      13'b0000001000000: n7774_o = 1'b0;
      13'b0000000100000: n7774_o = 1'b0;
      13'b0000000010000: n7774_o = 1'b0;
      13'b0000000001000: n7774_o = 1'b0;
      13'b0000000000100: n7774_o = 1'b0;
      13'b0000000000010: n7774_o = 1'b0;
      13'b0000000000001: n7774_o = n3135_o;
      default: n7774_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7776_o = 1'b0;
      13'b0100000000000: n7776_o = 1'b0;
      13'b0010000000000: n7776_o = 1'b0;
      13'b0001000000000: n7776_o = 1'b0;
      13'b0000100000000: n7776_o = 1'b0;
      13'b0000010000000: n7776_o = 1'b0;
      13'b0000001000000: n7776_o = 1'b0;
      13'b0000000100000: n7776_o = 1'b0;
      13'b0000000010000: n7776_o = 1'b0;
      13'b0000000001000: n7776_o = 1'b0;
      13'b0000000000100: n7776_o = n5847_o;
      13'b0000000000010: n7776_o = 1'b0;
      13'b0000000000001: n7776_o = 1'b0;
      default: n7776_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7778_o = 1'b0;
      13'b0100000000000: n7778_o = 1'b0;
      13'b0010000000000: n7778_o = 1'b0;
      13'b0001000000000: n7778_o = 1'b0;
      13'b0000100000000: n7778_o = 1'b0;
      13'b0000010000000: n7778_o = 1'b0;
      13'b0000001000000: n7778_o = 1'b0;
      13'b0000000100000: n7778_o = 1'b0;
      13'b0000000010000: n7778_o = 1'b0;
      13'b0000000001000: n7778_o = n6078_o;
      13'b0000000000100: n7778_o = 1'b0;
      13'b0000000000010: n7778_o = 1'b0;
      13'b0000000000001: n7778_o = 1'b0;
      default: n7778_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7780_o = 1'b0;
      13'b0100000000000: n7780_o = 1'b0;
      13'b0010000000000: n7780_o = n7079_o;
      13'b0001000000000: n7780_o = 1'b0;
      13'b0000100000000: n7780_o = 1'b0;
      13'b0000010000000: n7780_o = 1'b0;
      13'b0000001000000: n7780_o = 1'b0;
      13'b0000000100000: n7780_o = 1'b0;
      13'b0000000010000: n7780_o = 1'b0;
      13'b0000000001000: n7780_o = 1'b0;
      13'b0000000000100: n7780_o = 1'b0;
      13'b0000000000010: n7780_o = 1'b0;
      13'b0000000000001: n7780_o = 1'b0;
      default: n7780_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7782_o = 1'b0;
      13'b0100000000000: n7782_o = n7424_o;
      13'b0010000000000: n7782_o = 1'b0;
      13'b0001000000000: n7782_o = n6821_o;
      13'b0000100000000: n7782_o = 1'b0;
      13'b0000010000000: n7782_o = 1'b0;
      13'b0000001000000: n7782_o = n6486_o;
      13'b0000000100000: n7782_o = 1'b0;
      13'b0000000010000: n7782_o = 1'b0;
      13'b0000000001000: n7782_o = n6080_o;
      13'b0000000000100: n7782_o = n5849_o;
      13'b0000000000010: n7782_o = 1'b0;
      13'b0000000000001: n7782_o = n3137_o;
      default: n7782_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7784_o = 1'b0;
      13'b0100000000000: n7784_o = 1'b0;
      13'b0010000000000: n7784_o = 1'b0;
      13'b0001000000000: n7784_o = 1'b0;
      13'b0000100000000: n7784_o = 1'b0;
      13'b0000010000000: n7784_o = 1'b0;
      13'b0000001000000: n7784_o = 1'b0;
      13'b0000000100000: n7784_o = 1'b0;
      13'b0000000010000: n7784_o = 1'b0;
      13'b0000000001000: n7784_o = 1'b0;
      13'b0000000000100: n7784_o = n5851_o;
      13'b0000000000010: n7784_o = 1'b0;
      13'b0000000000001: n7784_o = 1'b0;
      default: n7784_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7786_o = 1'b0;
      13'b0100000000000: n7786_o = 1'b0;
      13'b0010000000000: n7786_o = 1'b0;
      13'b0001000000000: n7786_o = 1'b0;
      13'b0000100000000: n7786_o = 1'b0;
      13'b0000010000000: n7786_o = 1'b0;
      13'b0000001000000: n7786_o = 1'b0;
      13'b0000000100000: n7786_o = 1'b0;
      13'b0000000010000: n7786_o = 1'b0;
      13'b0000000001000: n7786_o = 1'b0;
      13'b0000000000100: n7786_o = n5853_o;
      13'b0000000000010: n7786_o = 1'b0;
      13'b0000000000001: n7786_o = 1'b0;
      default: n7786_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7788_o = 1'b0;
      13'b0100000000000: n7788_o = 1'b0;
      13'b0010000000000: n7788_o = 1'b0;
      13'b0001000000000: n7788_o = 1'b0;
      13'b0000100000000: n7788_o = 1'b0;
      13'b0000010000000: n7788_o = 1'b0;
      13'b0000001000000: n7788_o = 1'b0;
      13'b0000000100000: n7788_o = 1'b0;
      13'b0000000010000: n7788_o = 1'b0;
      13'b0000000001000: n7788_o = 1'b0;
      13'b0000000000100: n7788_o = n5855_o;
      13'b0000000000010: n7788_o = 1'b0;
      13'b0000000000001: n7788_o = 1'b0;
      default: n7788_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7790_o = 2'b00;
      13'b0100000000000: n7790_o = 2'b00;
      13'b0010000000000: n7790_o = 2'b00;
      13'b0001000000000: n7790_o = 2'b00;
      13'b0000100000000: n7790_o = 2'b00;
      13'b0000010000000: n7790_o = 2'b00;
      13'b0000001000000: n7790_o = 2'b00;
      13'b0000000100000: n7790_o = 2'b00;
      13'b0000000010000: n7790_o = 2'b00;
      13'b0000000001000: n7790_o = 2'b00;
      13'b0000000000100: n7790_o = n5858_o;
      13'b0000000000010: n7790_o = 2'b00;
      13'b0000000000001: n7790_o = 2'b00;
      default: n7790_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7792_o = 1'b0;
      13'b0100000000000: n7792_o = n7425_o;
      13'b0010000000000: n7792_o = n7081_o;
      13'b0001000000000: n7792_o = 1'b0;
      13'b0000100000000: n7792_o = 1'b0;
      13'b0000010000000: n7792_o = n6604_o;
      13'b0000001000000: n7792_o = n6487_o;
      13'b0000000100000: n7792_o = n6167_o;
      13'b0000000010000: n7792_o = 1'b0;
      13'b0000000001000: n7792_o = n6081_o;
      13'b0000000000100: n7792_o = n5860_o;
      13'b0000000000010: n7792_o = n3346_o;
      13'b0000000000001: n7792_o = n3138_o;
      default: n7792_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7794_o = 1'b0;
      13'b0100000000000: n7794_o = 1'b0;
      13'b0010000000000: n7794_o = n7083_o;
      13'b0001000000000: n7794_o = 1'b0;
      13'b0000100000000: n7794_o = 1'b0;
      13'b0000010000000: n7794_o = 1'b0;
      13'b0000001000000: n7794_o = 1'b0;
      13'b0000000100000: n7794_o = 1'b0;
      13'b0000000010000: n7794_o = 1'b0;
      13'b0000000001000: n7794_o = 1'b0;
      13'b0000000000100: n7794_o = 1'b0;
      13'b0000000000010: n7794_o = 1'b0;
      13'b0000000000001: n7794_o = 1'b0;
      default: n7794_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7796_o = 2'b00;
      13'b0100000000000: n7796_o = n7427_o;
      13'b0010000000000: n7796_o = 2'b00;
      13'b0001000000000: n7796_o = 2'b00;
      13'b0000100000000: n7796_o = 2'b00;
      13'b0000010000000: n7796_o = 2'b00;
      13'b0000001000000: n7796_o = 2'b00;
      13'b0000000100000: n7796_o = 2'b00;
      13'b0000000010000: n7796_o = 2'b00;
      13'b0000000001000: n7796_o = 2'b00;
      13'b0000000000100: n7796_o = 2'b00;
      13'b0000000000010: n7796_o = 2'b00;
      13'b0000000000001: n7796_o = 2'b00;
      default: n7796_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7798_o = 2'b00;
      13'b0100000000000: n7798_o = 2'b00;
      13'b0010000000000: n7798_o = 2'b00;
      13'b0001000000000: n7798_o = 2'b00;
      13'b0000100000000: n7798_o = 2'b00;
      13'b0000010000000: n7798_o = 2'b00;
      13'b0000001000000: n7798_o = n6489_o;
      13'b0000000100000: n7798_o = 2'b00;
      13'b0000000010000: n7798_o = 2'b00;
      13'b0000000001000: n7798_o = 2'b00;
      13'b0000000000100: n7798_o = 2'b00;
      13'b0000000000010: n7798_o = 2'b00;
      13'b0000000000001: n7798_o = 2'b00;
      default: n7798_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7800_o = 1'b0;
      13'b0100000000000: n7800_o = n7428_o;
      13'b0010000000000: n7800_o = 1'b0;
      13'b0001000000000: n7800_o = 1'b0;
      13'b0000100000000: n7800_o = 1'b0;
      13'b0000010000000: n7800_o = 1'b0;
      13'b0000001000000: n7800_o = 1'b0;
      13'b0000000100000: n7800_o = 1'b0;
      13'b0000000010000: n7800_o = 1'b0;
      13'b0000000001000: n7800_o = 1'b0;
      13'b0000000000100: n7800_o = 1'b0;
      13'b0000000000010: n7800_o = 1'b0;
      13'b0000000000001: n7800_o = 1'b0;
      default: n7800_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7802_o = 1'b0;
      13'b0100000000000: n7802_o = 1'b0;
      13'b0010000000000: n7802_o = 1'b0;
      13'b0001000000000: n7802_o = 1'b0;
      13'b0000100000000: n7802_o = 1'b0;
      13'b0000010000000: n7802_o = 1'b0;
      13'b0000001000000: n7802_o = 1'b0;
      13'b0000000100000: n7802_o = 1'b0;
      13'b0000000010000: n7802_o = 1'b0;
      13'b0000000001000: n7802_o = 1'b0;
      13'b0000000000100: n7802_o = n5861_o;
      13'b0000000000010: n7802_o = 1'b0;
      13'b0000000000001: n7802_o = 1'b0;
      default: n7802_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7573_o)
      13'b1000000000000: n7803_o = n2180_o;
      13'b0100000000000: n7803_o = n7429_o;
      13'b0010000000000: n7803_o = n2180_o;
      13'b0001000000000: n7803_o = n6822_o;
      13'b0000100000000: n7803_o = n2180_o;
      13'b0000010000000: n7803_o = n2180_o;
      13'b0000001000000: n7803_o = n6490_o;
      13'b0000000100000: n7803_o = n2180_o;
      13'b0000000010000: n7803_o = n6144_o;
      13'b0000000001000: n7803_o = n6082_o;
      13'b0000000000100: n7803_o = n5862_o;
      13'b0000000000010: n7803_o = n3313_o;
      13'b0000000000001: n7803_o = n3139_o;
      default: n7803_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7804_o = n2184_o ? make_berr : n7574_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7805_o = n2184_o ? n1921_o : n7576_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7806_o = n2184_o ? datatype : n7577_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7807_o = n2184_o ? n2026_o : n7578_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7808_o = n2184_o ? n2148_o : n7579_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7810_o = n2184_o ? 1'b0 : n7581_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7812_o = n2184_o ? n2151_o : n7582_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7814_o = n2184_o ? 1'b0 : n7584_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7817_o = n2184_o ? 1'b0 : n7586_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7819_o = n2184_o ? n2015_o : n7587_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7821_o = n2184_o ? 1'b0 : n7589_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7824_o = n2184_o ? 1'b0 : n7591_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7827_o = n2184_o ? 1'b0 : n7593_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7830_o = n2184_o ? 1'b0 : n7595_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7833_o = n2184_o ? 1'b0 : n7597_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7836_o = n2184_o ? 1'b0 : n7599_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7839_o = n2184_o ? 1'b0 : n7601_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7842_o = n2184_o ? 1'b0 : n7603_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7845_o = n2184_o ? 1'b0 : n7605_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7848_o = n2184_o ? 1'b0 : n7607_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7850_o = n2184_o ? n1900_o : n7608_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7851_o = n2184_o ? n1906_o : n7609_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7853_o = n2184_o ? 1'b0 : n7611_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7855_o = n2184_o ? n2154_o : n7612_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7857_o = n2184_o ? 1'b0 : n7615_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7861_o = n2184_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7864_o = n2184_o ? 1'b0 : n7617_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7867_o = n2184_o ? 1'b0 : n7620_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7870_o = n2184_o ? 1'b0 : n7622_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7873_o = n2184_o ? 1'b0 : n7624_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7876_o = n2184_o ? 1'b0 : n7626_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7879_o = n2184_o ? 1'b1 : n7631_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7882_o = n2184_o ? 1'b0 : n7633_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7885_o = n2184_o ? 1'b0 : n7635_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7888_o = n2184_o ? 1'b0 : n7637_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7891_o = n2184_o ? 1'b0 : n7639_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7894_o = n2184_o ? 1'b0 : n7641_o;
  assign n7896_o = {n7647_o, n7645_o};
  assign n7897_o = {n7664_o, n7662_o, n7660_o, n7659_o, n7657_o};
  assign n7898_o = {n7672_o, n7670_o, n7667_o};
  assign n7899_o = {n7712_o, n7710_o, n7708_o, n7705_o, n7701_o, n7698_o, n7695_o, n7692_o, n7690_o, n7687_o, n7684_o, n7678_o};
  assign n7900_o = {n7724_o, n7721_o};
  assign n7901_o = {n7734_o, n7732_o, n7730_o};
  assign n7902_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7903_o = n2184_o ? n7902_o : n7643_o;
  assign n7906_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7907_o = n2184_o ? n7906_o : n7649_o;
  assign n7908_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7909_o = n2184_o ? n7908_o : n7651_o;
  assign n7910_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7911_o = n2184_o ? n7910_o : n7653_o;
  assign n7912_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7913_o = n2184_o ? n7912_o : n7655_o;
  assign n7914_o = n1909_o[37:36];
  assign n7915_o = {n1940_o, n2007_o, n7914_o};
  assign n7917_o = n1909_o[44:42];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7918_o = n2184_o ? n7917_o : n7898_o;
  assign n7919_o = {n2179_o, n2168_o, n2177_o, n2166_o};
  assign n7921_o = n1909_o[67];
  assign n7922_o = {n7921_o, n2019_o, n2178_o};
  assign n7924_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7925_o = n2184_o ? n7924_o : n7717_o;
  assign n7926_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7927_o = n2184_o ? n7926_o : n7719_o;
  assign n7928_o = n1909_o[74];
  assign n7929_o = {n7928_o, n2171_o};
  assign n7931_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7932_o = n2184_o ? n7931_o : n7726_o;
  assign n7933_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7934_o = n2184_o ? n7933_o : n7728_o;
  assign n7938_o = n1909_o[21];
  assign n7939_o = n1909_o[16:1];
  assign n7940_o = n1909_o[23];
  assign n7945_o = n1909_o[33:30];
  assign n7946_o = n1909_o[35];
  assign n7947_o = n1909_o[45];
  assign n7950_o = n1909_o[68];
  assign n7951_o = n1909_o[72];
  assign n7952_o = n1909_o[70];
  assign n7956_o = n1909_o[81];
  assign n7958_o = {n7764_o, n7761_o, n7757_o, n7753_o, n7750_o, n7747_o, n7743_o, n7740_o, n7737_o};
  assign n7959_o = {n7778_o, n7776_o, n7774_o, n7772_o, n7770_o, n7768_o, n7766_o};
  assign n7960_o = {n7792_o, n7790_o, n7788_o, n7786_o};
  assign n7961_o = {n7798_o, n7796_o};
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7963_o = n2184_o ? 9'b000000000 : n7958_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7965_o = n2184_o ? 7'b0000000 : n7959_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7967_o = n2184_o ? 1'b0 : n7780_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7969_o = n2184_o ? 1'b0 : n7782_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7971_o = n2184_o ? 1'b0 : n7784_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7975_o = n2184_o ? 1'b0 : n7794_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7977_o = n2184_o ? 4'b0000 : n7961_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7979_o = n2184_o ? 1'b0 : n7800_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7981_o = n2184_o ? 1'b0 : n7802_o;
  assign n7985_o = n7982_o[9];
  assign n7987_o = n7982_o[19:17];
  assign n7991_o = n7982_o[27];
  assign n7993_o = n7982_o[29];
  assign n7995_o = n7982_o[66:35];
  assign n7997_o = n7982_o[74:68];
  assign n7999_o = n7982_o[80:79];
  assign n8000_o = n7982_o[87:82];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8001_o = n2184_o ? n2180_o : n7803_o;
  /* TG68KdotC_Kernel.vhd:3201:36  */
  assign n8002_o = set_exec[8];
  /* TG68KdotC_Kernel.vhd:3201:44  */
  assign n8003_o = ~n8002_o;
  /* TG68KdotC_Kernel.vhd:3201:60  */
  assign n8004_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:3201:63  */
  assign n8005_o = ~n8004_o;
  /* TG68KdotC_Kernel.vhd:3201:77  */
  assign n8006_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3201:89  */
  assign n8008_o = n8006_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3201:68  */
  assign n8009_o = n8005_o | n8008_o;
  /* TG68KdotC_Kernel.vhd:3201:49  */
  assign n8010_o = n8009_o & n8003_o;
  assign n8012_o = n7972_o[4];
  assign n8013_o = n7960_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8014_o = n2184_o ? n8012_o : n8013_o;
  /* TG68KdotC_Kernel.vhd:3201:25  */
  assign n8015_o = n8010_o ? 1'b1 : n8014_o;
  /* TG68KdotC_Kernel.vhd:3204:34  */
  assign n8016_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:3209:42  */
  assign n8018_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:3209:33  */
  assign n8020_o = n8018_o ? 1'b1 : n7830_o;
  /* TG68KdotC_Kernel.vhd:3212:33  */
  assign n8022_o = setexecopc ? 1'b1 : n7848_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8024_o = n8030_o ? 1'b1 : n7817_o;
  /* TG68KdotC_Kernel.vhd:3204:25  */
  assign n8025_o = n8016_o ? n7830_o : n8020_o;
  /* TG68KdotC_Kernel.vhd:3204:25  */
  assign n8027_o = n8016_o ? n7833_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3204:25  */
  assign n8028_o = n8016_o ? n7848_o : n8022_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8029_o = n8036_o ? 1'b1 : n7969_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8030_o = n8016_o & build_logical;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8031_o = build_logical ? n8025_o : n7830_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8032_o = build_logical ? n8027_o : n7833_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8033_o = build_logical ? n8028_o : n7848_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8035_o = build_logical ? 1'b1 : n7885_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8036_o = n8016_o & build_logical;
  assign n8037_o = n7972_o[4];
  assign n8038_o = n7960_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8039_o = n2184_o ? n8037_o : n8038_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n8040_o = build_logical ? n8015_o : n8039_o;
  assign n8041_o = n7972_o[3:0];
  assign n8042_o = n7960_o[3:0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8043_o = n2184_o ? n8041_o : n8042_o;
  /* TG68KdotC_Kernel.vhd:3224:34  */
  assign n8046_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:3226:50  */
  assign n8047_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:3226:62  */
  assign n8049_o = n8047_o == 3'b111;
  assign n8051_o = n7919_o[4];
  assign n8052_o = n7899_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8053_o = n2184_o ? n8051_o : n8052_o;
  /* TG68KdotC_Kernel.vhd:3226:41  */
  assign n8054_o = n8049_o ? 1'b1 : n8053_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8058_o = n8094_o ? 2'b10 : n7807_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8060_o = n8099_o ? 1'b1 : n7842_o;
  assign n8061_o = n7915_o[2];
  assign n8062_o = n7897_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8063_o = n2184_o ? n8061_o : n8062_o;
  /* TG68KdotC_Kernel.vhd:3225:33  */
  assign n8064_o = decodeopc ? 1'b1 : n8063_o;
  assign n8065_o = n7919_o[1];
  assign n8066_o = n7899_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8067_o = n2184_o ? n8065_o : n8066_o;
  /* TG68KdotC_Kernel.vhd:3225:33  */
  assign n8068_o = decodeopc ? 1'b1 : n8067_o;
  assign n8069_o = n7919_o[4];
  assign n8070_o = n7899_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8071_o = n2184_o ? n8069_o : n8070_o;
  /* TG68KdotC_Kernel.vhd:3225:33  */
  assign n8072_o = decodeopc ? n8054_o : n8071_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8074_o = n8134_o ? 7'b0100001 : n8001_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8076_o = decodeopc & n8046_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8077_o = decodeopc & n8046_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8079_o = n8046_o ? n8033_o : 1'b1;
  assign n8080_o = n7915_o[2];
  assign n8081_o = n7897_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8082_o = n2184_o ? n8080_o : n8081_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8083_o = n8046_o ? n8064_o : n8082_o;
  assign n8084_o = n7919_o[1];
  assign n8085_o = n7899_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8086_o = n2184_o ? n8084_o : n8085_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8087_o = n8046_o ? n8068_o : n8086_o;
  assign n8088_o = n7919_o[4];
  assign n8089_o = n7899_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8090_o = n2184_o ? n8088_o : n8089_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8091_o = n8046_o ? n8072_o : n8090_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8092_o = n8046_o ? n8040_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n8093_o = decodeopc & n8046_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8094_o = n8076_o & build_bcd;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8096_o = build_bcd ? 1'b1 : n8024_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8098_o = build_bcd ? 1'b1 : n8032_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8099_o = n8077_o & build_bcd;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8100_o = build_bcd ? n8079_o : n8033_o;
  assign n8101_o = n7915_o[2];
  assign n8102_o = n7897_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8103_o = n2184_o ? n8101_o : n8102_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8104_o = build_bcd ? n8083_o : n8103_o;
  assign n8105_o = n7919_o[1];
  assign n8106_o = n7899_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8107_o = n2184_o ? n8105_o : n8106_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8108_o = build_bcd ? n8087_o : n8107_o;
  assign n8109_o = n7919_o[4];
  assign n8110_o = n7899_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8111_o = n2184_o ? n8109_o : n8110_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8112_o = build_bcd ? n8091_o : n8111_o;
  assign n8122_o = n7919_o[0];
  assign n8123_o = n7899_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8124_o = n2184_o ? n8122_o : n8123_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8131_o = build_bcd ? 1'b1 : n8029_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8132_o = build_bcd ? 1'b1 : n7971_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8133_o = build_bcd ? n8092_o : n8040_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n8134_o = n8093_o & build_bcd;
  /* TG68KdotC_Kernel.vhd:3246:33  */
  assign n8135_o = ~trapd;
  /* TG68KdotC_Kernel.vhd:3244:17  */
  assign n8137_o = n8138_o ? 1'b1 : n7821_o;
  /* TG68KdotC_Kernel.vhd:3244:17  */
  assign n8138_o = n8135_o & set_z_error;
  /* TG68KdotC_Kernel.vhd:3244:17  */
  assign n8140_o = set_z_error ? 1'b1 : n7879_o;
  /* TG68KdotC_Kernel.vhd:3257:25  */
  assign n8142_o = clkena_lw ? trapmake : trapd;
  /* TG68KdotC_Kernel.vhd:3257:25  */
  assign n8143_o = clkena_lw ? next_micro_state : micro_state;
  /* TG68KdotC_Kernel.vhd:3255:17  */
  assign n8144_o = reset ? trapd : n8142_o;
  /* TG68KdotC_Kernel.vhd:3255:17  */
  assign n8146_o = reset ? 7'b0000010 : n8143_o;
  /* TG68KdotC_Kernel.vhd:3264:33  */
  assign n8152_o = micro_state == 7'b0000010;
  /* TG68KdotC_Kernel.vhd:3269:33  */
  assign n8155_o = micro_state == 7'b0000011;
  /* TG68KdotC_Kernel.vhd:3274:33  */
  assign n8158_o = micro_state == 7'b0000100;
  /* TG68KdotC_Kernel.vhd:3280:49  */
  assign n8159_o = brief[8];
  /* TG68KdotC_Kernel.vhd:3280:52  */
  assign n8160_o = ~n8159_o;
  /* TG68KdotC_Kernel.vhd:3280:57  */
  assign n8162_o = n8160_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3280:82  */
  assign n8163_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3280:85  */
  assign n8164_o = ~n8163_o;
  /* TG68KdotC_Kernel.vhd:3280:90  */
  assign n8166_o = 1'b1 & n8164_o;
  /* TG68KdotC_Kernel.vhd:3280:75  */
  assign n8167_o = n8162_o | n8166_o;
  /* TG68KdotC_Kernel.vhd:3287:57  */
  assign n8169_o = brief[7];
  /* TG68KdotC_Kernel.vhd:3289:59  */
  assign n8170_o = exec[22];
  /* TG68KdotC_Kernel.vhd:3289:49  */
  assign n8172_o = n8170_o ? 1'b1 : n2164_o;
  /* TG68KdotC_Kernel.vhd:3287:49  */
  assign n8174_o = n8169_o ? 1'b1 : n2157_o;
  /* TG68KdotC_Kernel.vhd:3287:49  */
  assign n8175_o = n8169_o ? n2164_o : n8172_o;
  /* TG68KdotC_Kernel.vhd:3292:57  */
  assign n8176_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3292:60  */
  assign n8177_o = ~n8176_o;
  /* TG68KdotC_Kernel.vhd:3295:65  */
  assign n8178_o = brief[4];
  assign n8180_o = n7929_o[0];
  assign n8181_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8182_o = n2184_o ? n8180_o : n8181_o;
  /* TG68KdotC_Kernel.vhd:3295:57  */
  assign n8183_o = n8178_o ? 1'b1 : n8182_o;
  /* TG68KdotC_Kernel.vhd:3292:49  */
  assign n8185_o = n8177_o ? 2'b01 : n8058_o;
  assign n8186_o = n7929_o[0];
  assign n8187_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8188_o = n2184_o ? n8186_o : n8187_o;
  /* TG68KdotC_Kernel.vhd:3292:49  */
  assign n8189_o = n8177_o ? n8188_o : n8183_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8191_o = n8167_o ? 2'b01 : n8185_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8194_o = n8167_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8197_o = n8167_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8198_o = n8167_o ? n2157_o : n8174_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8199_o = n8167_o ? n2164_o : n8175_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8200_o = n8167_o ? 1'b1 : n7952_o;
  assign n8201_o = n7929_o[0];
  assign n8202_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8203_o = n2184_o ? n8201_o : n8202_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8204_o = n8167_o ? n8203_o : n8189_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8207_o = n8167_o ? 7'b0000110 : 7'b0001011;
  /* TG68KdotC_Kernel.vhd:3279:33  */
  assign n8209_o = micro_state == 7'b0000101;
  /* TG68KdotC_Kernel.vhd:3302:33  */
  assign n8212_o = micro_state == 7'b0000110;
  /* TG68KdotC_Kernel.vhd:3310:49  */
  assign n8213_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3310:41  */
  assign n8216_o = n8213_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3313:49  */
  assign n8217_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3313:52  */
  assign n8218_o = ~n8217_o;
  /* TG68KdotC_Kernel.vhd:3313:66  */
  assign n8219_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3313:69  */
  assign n8220_o = ~n8219_o;
  /* TG68KdotC_Kernel.vhd:3313:57  */
  assign n8221_o = n8220_o & n8218_o;
  /* TG68KdotC_Kernel.vhd:3316:57  */
  assign n8223_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3316:69  */
  assign n8225_o = n8223_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3316:49  */
  assign n8228_o = n8225_o ? 7'b0000110 : 7'b0001100;
  /* TG68KdotC_Kernel.vhd:3322:57  */
  assign n8229_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3322:69  */
  assign n8231_o = n8229_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8235_o = n8231_o ? n8058_o : 2'b10;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8238_o = n8231_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8240_o = n8231_o ? 1'b1 : n7808_o;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8241_o = n8231_o ? 1'b1 : n2170_o;
  assign n8242_o = n7929_o[0];
  assign n8243_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8244_o = n2184_o ? n8242_o : n8243_o;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8245_o = n8231_o ? n8244_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8247_o = n8231_o ? n8074_o : 7'b0001101;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8249_o = n8221_o ? 2'b01 : n8235_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8251_o = n8221_o ? 1'b0 : n8238_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8252_o = n8221_o ? n7808_o : n8240_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8253_o = n8221_o ? n2170_o : n8241_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8254_o = n8221_o ? 1'b1 : n7952_o;
  assign n8255_o = n7929_o[0];
  assign n8256_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8257_o = n2184_o ? n8255_o : n8256_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8258_o = n8221_o ? n8257_o : n8245_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8259_o = n8221_o ? n8228_o : n8247_o;
  /* TG68KdotC_Kernel.vhd:3309:33  */
  assign n8261_o = micro_state == 7'b0001011;
  /* TG68KdotC_Kernel.vhd:3333:33  */
  assign n8264_o = micro_state == 7'b0001100;
  /* TG68KdotC_Kernel.vhd:3343:49  */
  assign n8266_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3343:52  */
  assign n8267_o = ~n8266_o;
  /* TG68KdotC_Kernel.vhd:3346:57  */
  assign n8268_o = brief[0];
  assign n8270_o = n7929_o[0];
  assign n8271_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8272_o = n2184_o ? n8270_o : n8271_o;
  /* TG68KdotC_Kernel.vhd:3346:49  */
  assign n8273_o = n8268_o ? 1'b1 : n8272_o;
  /* TG68KdotC_Kernel.vhd:3343:41  */
  assign n8275_o = n8267_o ? 2'b01 : n8058_o;
  assign n8276_o = n7929_o[0];
  assign n8277_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8278_o = n2184_o ? n8276_o : n8277_o;
  /* TG68KdotC_Kernel.vhd:3343:41  */
  assign n8279_o = n8267_o ? n8278_o : n8273_o;
  /* TG68KdotC_Kernel.vhd:3340:33  */
  assign n8281_o = micro_state == 7'b0001101;
  /* TG68KdotC_Kernel.vhd:3353:49  */
  assign n8282_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3353:41  */
  assign n8285_o = n8282_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3356:49  */
  assign n8286_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3356:52  */
  assign n8287_o = ~n8286_o;
  /* TG68KdotC_Kernel.vhd:3356:66  */
  assign n8288_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3356:57  */
  assign n8289_o = n8288_o & n8287_o;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8293_o = n8289_o ? 2'b01 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8295_o = n8289_o ? n7808_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8296_o = n8289_o ? n2170_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8297_o = n8289_o ? 1'b1 : n7952_o;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8299_o = n8289_o ? 7'b0000110 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3352:33  */
  assign n8301_o = micro_state == 7'b0001110;
  /* TG68KdotC_Kernel.vhd:3366:33  */
  assign n8303_o = micro_state == 7'b0000111;
  /* TG68KdotC_Kernel.vhd:3372:49  */
  assign n8304_o = brief[8];
  /* TG68KdotC_Kernel.vhd:3372:52  */
  assign n8305_o = ~n8304_o;
  /* TG68KdotC_Kernel.vhd:3372:57  */
  assign n8307_o = n8305_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3372:82  */
  assign n8308_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3372:85  */
  assign n8309_o = ~n8308_o;
  /* TG68KdotC_Kernel.vhd:3372:90  */
  assign n8311_o = 1'b1 & n8309_o;
  /* TG68KdotC_Kernel.vhd:3372:75  */
  assign n8312_o = n8307_o | n8311_o;
  /* TG68KdotC_Kernel.vhd:3379:57  */
  assign n8314_o = brief[7];
  /* TG68KdotC_Kernel.vhd:3379:49  */
  assign n8316_o = n8314_o ? 1'b1 : n2157_o;
  /* TG68KdotC_Kernel.vhd:3384:57  */
  assign n8317_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3384:60  */
  assign n8318_o = ~n8317_o;
  /* TG68KdotC_Kernel.vhd:3387:65  */
  assign n8319_o = brief[4];
  assign n8321_o = n7929_o[0];
  assign n8322_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8323_o = n2184_o ? n8321_o : n8322_o;
  /* TG68KdotC_Kernel.vhd:3387:57  */
  assign n8324_o = n8319_o ? 1'b1 : n8323_o;
  /* TG68KdotC_Kernel.vhd:3384:49  */
  assign n8326_o = n8318_o ? 2'b01 : n8058_o;
  assign n8327_o = n7929_o[0];
  assign n8328_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8329_o = n2184_o ? n8327_o : n8328_o;
  /* TG68KdotC_Kernel.vhd:3384:49  */
  assign n8330_o = n8318_o ? n8329_o : n8324_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8332_o = n8312_o ? 2'b01 : n8326_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8335_o = n8312_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8338_o = n8312_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8339_o = n8312_o ? n2157_o : n8316_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8340_o = n8312_o ? 1'b1 : n7952_o;
  assign n8341_o = n7929_o[0];
  assign n8342_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8343_o = n2184_o ? n8341_o : n8342_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8344_o = n8312_o ? n8343_o : n8330_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8347_o = n8312_o ? 7'b0010100 : 7'b0001111;
  /* TG68KdotC_Kernel.vhd:3371:33  */
  assign n8349_o = micro_state == 7'b0010011;
  /* TG68KdotC_Kernel.vhd:3394:33  */
  assign n8352_o = micro_state == 7'b0010100;
  /* TG68KdotC_Kernel.vhd:3403:49  */
  assign n8353_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3403:41  */
  assign n8356_o = n8353_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3406:49  */
  assign n8357_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3406:52  */
  assign n8358_o = ~n8357_o;
  /* TG68KdotC_Kernel.vhd:3406:66  */
  assign n8359_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3406:69  */
  assign n8360_o = ~n8359_o;
  /* TG68KdotC_Kernel.vhd:3406:57  */
  assign n8361_o = n8360_o & n8358_o;
  /* TG68KdotC_Kernel.vhd:3409:57  */
  assign n8363_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3409:69  */
  assign n8365_o = n8363_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3409:49  */
  assign n8368_o = n8365_o ? 7'b0010100 : 7'b0010000;
  /* TG68KdotC_Kernel.vhd:3415:57  */
  assign n8369_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3415:69  */
  assign n8371_o = n8369_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8376_o = n8371_o ? 2'b11 : 2'b10;
  assign n8377_o = n7922_o[1];
  assign n8378_o = n7715_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8379_o = n2184_o ? n8377_o : n8378_o;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8380_o = n8371_o ? n8379_o : 1'b1;
  assign n8381_o = n7929_o[0];
  assign n8382_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8383_o = n2184_o ? n8381_o : n8382_o;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8384_o = n8371_o ? n8383_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8387_o = n8371_o ? 7'b0000001 : 7'b0010001;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8389_o = n8361_o ? 2'b01 : n8376_o;
  assign n8390_o = n7922_o[1];
  assign n8391_o = n7715_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8392_o = n2184_o ? n8390_o : n8391_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8393_o = n8361_o ? n8392_o : n8380_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8394_o = n8361_o ? 1'b1 : n7952_o;
  assign n8395_o = n7929_o[0];
  assign n8396_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8397_o = n2184_o ? n8395_o : n8396_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8398_o = n8361_o ? n8397_o : n8384_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8399_o = n8361_o ? n8368_o : n8387_o;
  /* TG68KdotC_Kernel.vhd:3402:33  */
  assign n8401_o = micro_state == 7'b0001111;
  /* TG68KdotC_Kernel.vhd:3426:33  */
  assign n8405_o = micro_state == 7'b0010000;
  /* TG68KdotC_Kernel.vhd:3437:49  */
  assign n8408_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3437:52  */
  assign n8409_o = ~n8408_o;
  /* TG68KdotC_Kernel.vhd:3440:57  */
  assign n8410_o = brief[0];
  assign n8412_o = n7929_o[0];
  assign n8413_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8414_o = n2184_o ? n8412_o : n8413_o;
  /* TG68KdotC_Kernel.vhd:3440:49  */
  assign n8415_o = n8410_o ? 1'b1 : n8414_o;
  /* TG68KdotC_Kernel.vhd:3437:41  */
  assign n8417_o = n8409_o ? 2'b01 : n8058_o;
  assign n8418_o = n7929_o[0];
  assign n8419_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8420_o = n2184_o ? n8418_o : n8419_o;
  /* TG68KdotC_Kernel.vhd:3437:41  */
  assign n8421_o = n8409_o ? n8420_o : n8415_o;
  /* TG68KdotC_Kernel.vhd:3433:33  */
  assign n8423_o = micro_state == 7'b0010001;
  /* TG68KdotC_Kernel.vhd:3448:49  */
  assign n8425_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3448:41  */
  assign n8428_o = n8425_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3451:49  */
  assign n8429_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3451:52  */
  assign n8430_o = ~n8429_o;
  /* TG68KdotC_Kernel.vhd:3451:66  */
  assign n8431_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3451:57  */
  assign n8432_o = n8431_o & n8430_o;
  /* TG68KdotC_Kernel.vhd:3451:41  */
  assign n8436_o = n8432_o ? 2'b01 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3451:41  */
  assign n8437_o = n8432_o ? 1'b1 : n7952_o;
  /* TG68KdotC_Kernel.vhd:3451:41  */
  assign n8440_o = n8432_o ? 7'b0010100 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3446:33  */
  assign n8442_o = micro_state == 7'b0010010;
  /* TG68KdotC_Kernel.vhd:3462:41  */
  assign n8444_o = exe_condition ? 1'b1 : n7804_o;
  /* TG68KdotC_Kernel.vhd:3462:41  */
  assign n8447_o = exe_condition ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3462:41  */
  assign n8449_o = exe_condition ? 7'b0000001 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3461:33  */
  assign n8451_o = micro_state == 7'b0010101;
  /* TG68KdotC_Kernel.vhd:3468:33  */
  assign n8453_o = micro_state == 7'b0010110;
  /* TG68KdotC_Kernel.vhd:3473:54  */
  assign n8454_o = ~long_start;
  /* TG68KdotC_Kernel.vhd:3473:41  */
  assign n8457_o = n8454_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3472:33  */
  assign n8460_o = micro_state == 7'b0010111;
  /* TG68KdotC_Kernel.vhd:3482:33  */
  assign n8462_o = micro_state == 7'b0011000;
  /* TG68KdotC_Kernel.vhd:3486:57  */
  assign n8463_o = ~exe_condition;
  /* TG68KdotC_Kernel.vhd:3488:57  */
  assign n8464_o = c_out[1];
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8466_o = n8472_o ? 1'b1 : n7804_o;
  /* TG68KdotC_Kernel.vhd:3488:49  */
  assign n8469_o = n8464_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8471_o = n8478_o ? 7'b0000001 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8472_o = n8464_o & n8463_o;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8475_o = n8463_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8477_o = n8463_o ? n8469_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8478_o = n8464_o & n8463_o;
  /* TG68KdotC_Kernel.vhd:3485:33  */
  assign n8480_o = micro_state == 7'b0011001;
  /* TG68KdotC_Kernel.vhd:3495:33  */
  assign n8486_o = micro_state == 7'b1000001;
  /* TG68KdotC_Kernel.vhd:3504:50  */
  assign n8487_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3507:58  */
  assign n8488_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3507:71  */
  assign n8490_o = n8488_o == 2'b00;
  assign n8492_o = n1909_o[88];
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8493_o = n8500_o ? 1'b1 : n8492_o;
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8495_o = n8487_o ? 2'b10 : n7806_o;
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8498_o = n8487_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8500_o = n8490_o & n8487_o;
  /* TG68KdotC_Kernel.vhd:3502:33  */
  assign n8505_o = micro_state == 7'b1000010;
  /* TG68KdotC_Kernel.vhd:3519:50  */
  assign n8507_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3519:41  */
  assign n8509_o = n8507_o ? 2'b10 : n7806_o;
  /* TG68KdotC_Kernel.vhd:3519:41  */
  assign n8512_o = n8507_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3526:61  */
  assign n8516_o = exec[88];
  /* TG68KdotC_Kernel.vhd:3527:50  */
  assign n8517_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:3527:41  */
  assign n8519_o = n8517_o ? 2'b01 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3527:41  */
  assign n8521_o = n8517_o ? 7'b1000100 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3516:33  */
  assign n8523_o = micro_state == 7'b1000011;
  /* TG68KdotC_Kernel.vhd:3531:33  */
  assign n8525_o = micro_state == 7'b1000100;
  /* TG68KdotC_Kernel.vhd:3535:49  */
  assign n8526_o = flags[0];
  /* TG68KdotC_Kernel.vhd:3535:41  */
  assign n8528_o = n8526_o ? 1'b1 : n8140_o;
  /* TG68KdotC_Kernel.vhd:3534:33  */
  assign n8530_o = micro_state == 7'b1000101;
  /* TG68KdotC_Kernel.vhd:3540:33  */
  assign n8532_o = micro_state == 7'b0110111;
  /* TG68KdotC_Kernel.vhd:3545:49  */
  assign n8533_o = flags[2];
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8540_o = n8533_o ? 2'b11 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8543_o = n8533_o ? 1'b0 : 1'b1;
  assign n8544_o = n1909_o[27];
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8545_o = n8533_o ? n8544_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8546_o = n8533_o ? n7913_o : 1'b1;
  assign n8547_o = n7915_o[4];
  assign n8548_o = n7897_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8549_o = n2184_o ? n8547_o : n8548_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8550_o = n8533_o ? 1'b1 : n8549_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8551_o = n8533_o ? 1'b1 : n1925_o;
  assign n8552_o = n1909_o[85];
  assign n8553_o = n7901_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8554_o = n2184_o ? n8552_o : n8553_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8555_o = n8533_o ? n8554_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8557_o = n8533_o ? 7'b0000001 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3543:33  */
  assign n8559_o = micro_state == 7'b0111000;
  /* TG68KdotC_Kernel.vhd:3559:63  */
  assign n8560_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3557:33  */
  assign n8563_o = micro_state == 7'b0111001;
  /* TG68KdotC_Kernel.vhd:3562:33  */
  assign n8569_o = micro_state == 7'b0111010;
  /* TG68KdotC_Kernel.vhd:3570:33  */
  assign n8572_o = micro_state == 7'b0111011;
  /* TG68KdotC_Kernel.vhd:3575:49  */
  assign n8573_o = flags[2];
  assign n8575_o = n1909_o[86];
  assign n8576_o = n7901_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8577_o = n2184_o ? n8575_o : n8576_o;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8578_o = n8573_o ? 1'b1 : n8577_o;
  /* TG68KdotC_Kernel.vhd:3574:33  */
  assign n8584_o = micro_state == 7'b0111100;
  /* TG68KdotC_Kernel.vhd:3585:33  */
  assign n8587_o = micro_state == 7'b0111101;
  /* TG68KdotC_Kernel.vhd:3590:49  */
  assign n8588_o = flags[2];
  /* TG68KdotC_Kernel.vhd:3594:71  */
  assign n8590_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8598_o = n8588_o ? 2'b11 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8601_o = n8588_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8603_o = n8588_o ? n8590_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8606_o = n8588_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8608_o = n8588_o ? 1'b1 : n7845_o;
  assign n8609_o = n1909_o[27];
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8610_o = n8588_o ? n8609_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8611_o = n8588_o ? n7913_o : 1'b1;
  assign n8612_o = n7915_o[4];
  assign n8613_o = n7897_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8614_o = n2184_o ? n8612_o : n8613_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8615_o = n8588_o ? 1'b1 : n8614_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8616_o = n8588_o ? 1'b1 : n2170_o;
  assign n8617_o = n7922_o[1];
  assign n8618_o = n7715_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8619_o = n2184_o ? n8617_o : n8618_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8620_o = n8588_o ? n8619_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8621_o = n8588_o ? n7934_o : 1'b1;
  assign n8622_o = n1909_o[85];
  assign n8623_o = n7901_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8624_o = n2184_o ? n8622_o : n8623_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8625_o = n8588_o ? n8624_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8628_o = n8588_o ? 7'b0111111 : 7'b1000000;
  /* TG68KdotC_Kernel.vhd:3589:33  */
  assign n8630_o = micro_state == 7'b0111110;
  /* TG68KdotC_Kernel.vhd:3607:33  */
  assign n8634_o = micro_state == 7'b0111111;
  /* TG68KdotC_Kernel.vhd:3614:33  */
  assign n8638_o = micro_state == 7'b1000000;
  /* TG68KdotC_Kernel.vhd:3620:58  */
  assign n8639_o = last_data_read[15:0];
  /* TG68KdotC_Kernel.vhd:3620:71  */
  assign n8641_o = n8639_o != 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3622:58  */
  assign n8642_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3622:70  */
  assign n8644_o = n8642_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3624:63  */
  assign n8646_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8648_o = n8656_o ? 1'b1 : n7913_o;
  /* TG68KdotC_Kernel.vhd:3622:49  */
  assign n8649_o = n8646_o & n8644_o;
  assign n8650_o = n7919_o[9];
  assign n8651_o = n7899_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8652_o = n2184_o ? n8650_o : n8651_o;
  /* TG68KdotC_Kernel.vhd:3622:49  */
  assign n8653_o = n8644_o ? 1'b1 : n8652_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8655_o = n8641_o ? 2'b01 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8656_o = n8649_o & n8641_o;
  assign n8657_o = n7919_o[9];
  assign n8658_o = n7899_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8659_o = n2184_o ? n8657_o : n8658_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8660_o = n8641_o ? n8653_o : n8659_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8662_o = n8641_o ? 7'b0011011 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3619:33  */
  assign n8664_o = micro_state == 7'b0011010;
  /* TG68KdotC_Kernel.vhd:3631:53  */
  assign n8665_o = ~movem_run;
  /* TG68KdotC_Kernel.vhd:3637:58  */
  assign n8668_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:3637:62  */
  assign n8669_o = ~n8668_o;
  /* TG68KdotC_Kernel.vhd:3637:49  */
  assign n8673_o = n8669_o ? 2'b11 : 2'b10;
  assign n8674_o = n7915_o[4];
  assign n8675_o = n7897_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8676_o = n2184_o ? n8674_o : n8675_o;
  /* TG68KdotC_Kernel.vhd:3637:49  */
  assign n8677_o = n8669_o ? 1'b1 : n8676_o;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8679_o = n8665_o ? 2'b01 : n8673_o;
  assign n8680_o = n7915_o[4];
  assign n8681_o = n7897_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8682_o = n2184_o ? n8680_o : n8681_o;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8683_o = n8665_o ? n8682_o : n8677_o;
  assign n8684_o = n7919_o[9];
  assign n8685_o = n7899_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8686_o = n2184_o ? n8684_o : n8685_o;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8687_o = n8665_o ? n8686_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8688_o = n8665_o ? n7925_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8690_o = n8665_o ? n8074_o : 7'b0011011;
  /* TG68KdotC_Kernel.vhd:3630:33  */
  assign n8692_o = micro_state == 7'b0011011;
  /* TG68KdotC_Kernel.vhd:3646:50  */
  assign n8693_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3646:62  */
  assign n8695_o = n8693_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3646:41  */
  assign n8697_o = n8695_o ? 1'b1 : n7808_o;
  /* TG68KdotC_Kernel.vhd:3645:33  */
  assign n8699_o = micro_state == 7'b0011101;
  /* TG68KdotC_Kernel.vhd:3651:50  */
  assign n8700_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:3651:62  */
  assign n8702_o = n8700_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3651:41  */
  assign n8704_o = n8702_o ? 1'b1 : n8112_o;
  /* TG68KdotC_Kernel.vhd:3650:33  */
  assign n8709_o = micro_state == 7'b0011110;
  /* TG68KdotC_Kernel.vhd:3661:50  */
  assign n8710_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3661:63  */
  assign n8712_o = n8710_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3661:41  */
  assign n8714_o = n8712_o ? 1'b1 : n8112_o;
  /* TG68KdotC_Kernel.vhd:3666:50  */
  assign n8716_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:3666:63  */
  assign n8718_o = n8716_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:3666:41  */
  assign n8721_o = n8718_o ? 2'b00 : 2'b01;
  /* TG68KdotC_Kernel.vhd:3660:33  */
  assign n8724_o = micro_state == 7'b0011111;
  /* TG68KdotC_Kernel.vhd:3676:33  */
  assign n8726_o = micro_state == 7'b0100000;
  /* TG68KdotC_Kernel.vhd:3680:50  */
  assign n8727_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3680:63  */
  assign n8729_o = n8727_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3680:41  */
  assign n8731_o = n8729_o ? 1'b1 : n8112_o;
  /* TG68KdotC_Kernel.vhd:3679:33  */
  assign n8734_o = micro_state == 7'b0100001;
  /* TG68KdotC_Kernel.vhd:3690:50  */
  assign n8735_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3690:63  */
  assign n8737_o = n8735_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3690:41  */
  assign n8739_o = n8737_o ? 1'b1 : n8112_o;
  /* TG68KdotC_Kernel.vhd:3689:33  */
  assign n8742_o = micro_state == 7'b0100010;
  /* TG68KdotC_Kernel.vhd:3699:33  */
  assign n8746_o = micro_state == 7'b0100011;
  /* TG68KdotC_Kernel.vhd:3705:33  */
  assign n8749_o = micro_state == 7'b0100100;
  /* TG68KdotC_Kernel.vhd:3709:33  */
  assign n8752_o = micro_state == 7'b0100101;
  /* TG68KdotC_Kernel.vhd:3714:33  */
  assign n8755_o = micro_state == 7'b0100110;
  /* TG68KdotC_Kernel.vhd:3718:33  */
  assign n8758_o = micro_state == 7'b0110010;
  /* TG68KdotC_Kernel.vhd:3735:71  */
  assign n8761_o = trap_interrupt | trap_trace;
  /* TG68KdotC_Kernel.vhd:3735:89  */
  assign n8762_o = n8761_o | trap_berr;
  /* TG68KdotC_Kernel.vhd:3735:49  */
  assign n8764_o = n8762_o ? 1'b1 : n8137_o;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8767_o = use_vbr_stackframe ? 2'b01 : 2'b10;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8768_o = use_vbr_stackframe ? n8137_o : n8764_o;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8769_o = use_vbr_stackframe ? 1'b1 : n1960_o;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8772_o = use_vbr_stackframe ? 7'b0110100 : 7'b0110101;
  /* TG68KdotC_Kernel.vhd:3725:33  */
  assign n8774_o = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:3743:63  */
  assign n8775_o = trap_interrupt | trap_trace;
  /* TG68KdotC_Kernel.vhd:3743:41  */
  assign n8777_o = n8775_o ? 1'b1 : n8137_o;
  /* TG68KdotC_Kernel.vhd:3742:33  */
  assign n8780_o = micro_state == 7'b0110100;
  /* TG68KdotC_Kernel.vhd:3751:33  */
  assign n8783_o = micro_state == 7'b0110101;
  /* TG68KdotC_Kernel.vhd:3758:33  */
  assign n8787_o = micro_state == 7'b0110110;
  /* TG68KdotC_Kernel.vhd:3770:33  */
  assign n8790_o = micro_state == 7'b1000110;
  /* TG68KdotC_Kernel.vhd:3776:33  */
  assign n8793_o = micro_state == 7'b1000111;
  /* TG68KdotC_Kernel.vhd:3782:33  */
  assign n8796_o = micro_state == 7'b1001000;
  /* TG68KdotC_Kernel.vhd:3788:33  */
  assign n8799_o = micro_state == 7'b1011011;
  /* TG68KdotC_Kernel.vhd:3794:33  */
  assign n8802_o = micro_state == 7'b1011100;
  /* TG68KdotC_Kernel.vhd:3800:33  */
  assign n8805_o = micro_state == 7'b1011101;
  /* TG68KdotC_Kernel.vhd:3806:33  */
  assign n8808_o = micro_state == 7'b1011110;
  /* TG68KdotC_Kernel.vhd:3826:62  */
  assign n8811_o = ~use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:3826:76  */
  assign n8812_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:3826:67  */
  assign n8813_o = n8811_o | n8812_o;
  /* TG68KdotC_Kernel.vhd:3826:41  */
  assign n8816_o = n8813_o ? 1'b1 : n7946_o;
  assign n8817_o = n7919_o[12];
  assign n8818_o = n7899_o[12];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8819_o = n2184_o ? n8817_o : n8818_o;
  /* TG68KdotC_Kernel.vhd:3826:41  */
  assign n8820_o = n8813_o ? 1'b1 : n8819_o;
  /* TG68KdotC_Kernel.vhd:3820:33  */
  assign n8822_o = micro_state == 7'b0101011;
  /* TG68KdotC_Kernel.vhd:3834:77  */
  assign n8824_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:3834:80  */
  assign n8825_o = ~n8824_o;
  /* TG68KdotC_Kernel.vhd:3834:67  */
  assign n8826_o = n8825_o & use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8829_o = n8826_o ? 2'b10 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8831_o = n8826_o ? 1'b1 : n7819_o;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8832_o = n8826_o ? 1'b1 : n8124_o;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8835_o = n8826_o ? 7'b0101101 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3831:33  */
  assign n8837_o = micro_state == 7'b0101100;
  /* TG68KdotC_Kernel.vhd:3847:33  */
  assign n8839_o = micro_state == 7'b0101101;
  /* TG68KdotC_Kernel.vhd:3854:56  */
  assign n8840_o = last_data_in[15:12];
  /* TG68KdotC_Kernel.vhd:3854:70  */
  assign n8842_o = n8840_o == 4'b0010;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8846_o = n8842_o ? 2'b10 : 2'b01;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8848_o = n8842_o ? 2'b10 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8850_o = n8842_o ? 1'b1 : n7819_o;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8851_o = n8842_o ? 1'b1 : n8124_o;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8854_o = n8842_o ? 7'b0101111 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3852:33  */
  assign n8856_o = micro_state == 7'b0101110;
  /* TG68KdotC_Kernel.vhd:3865:33  */
  assign n8858_o = micro_state == 7'b0101111;
  /* TG68KdotC_Kernel.vhd:3869:33  */
  assign n8860_o = micro_state == 7'b0110000;
  /* TG68KdotC_Kernel.vhd:3871:33  */
  assign n8863_o = micro_state == 7'b0110001;
  /* TG68KdotC_Kernel.vhd:3878:50  */
  assign n8865_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:63  */
  assign n8867_o = n8865_o == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:3878:79  */
  assign n8868_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:92  */
  assign n8870_o = n8868_o == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:3878:71  */
  assign n8871_o = n8867_o | n8870_o;
  /* TG68KdotC_Kernel.vhd:3878:108  */
  assign n8872_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:121  */
  assign n8874_o = n8872_o == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:3878:100  */
  assign n8875_o = n8871_o | n8874_o;
  /* TG68KdotC_Kernel.vhd:3878:137  */
  assign n8876_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:150  */
  assign n8878_o = n8876_o == 12'b100000000001;
  /* TG68KdotC_Kernel.vhd:3878:129  */
  assign n8879_o = n8875_o | n8878_o;
  /* TG68KdotC_Kernel.vhd:3879:48  */
  assign n8880_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3879:66  */
  assign n8881_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:79  */
  assign n8883_o = n8881_o == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:3879:95  */
  assign n8884_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:108  */
  assign n8886_o = n8884_o == 12'b100000000010;
  /* TG68KdotC_Kernel.vhd:3879:87  */
  assign n8887_o = n8883_o | n8886_o;
  /* TG68KdotC_Kernel.vhd:3879:124  */
  assign n8888_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:137  */
  assign n8890_o = n8888_o == 12'b100000000011;
  /* TG68KdotC_Kernel.vhd:3879:116  */
  assign n8891_o = n8887_o | n8890_o;
  /* TG68KdotC_Kernel.vhd:3879:153  */
  assign n8892_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:166  */
  assign n8894_o = n8892_o == 12'b100000000100;
  /* TG68KdotC_Kernel.vhd:3879:145  */
  assign n8895_o = n8891_o | n8894_o;
  /* TG68KdotC_Kernel.vhd:3879:56  */
  assign n8896_o = n8895_o & n8880_o;
  /* TG68KdotC_Kernel.vhd:3878:159  */
  assign n8897_o = n8879_o | n8896_o;
  /* TG68KdotC_Kernel.vhd:3880:58  */
  assign n8898_o = opcode[0];
  /* TG68KdotC_Kernel.vhd:3880:61  */
  assign n8899_o = ~n8898_o;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8901_o = n8906_o ? 1'b1 : n7913_o;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8903_o = n8897_o ? n7857_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8905_o = n8897_o ? n8140_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8906_o = n8899_o & n8897_o;
  /* TG68KdotC_Kernel.vhd:3875:33  */
  assign n8908_o = micro_state == 7'b1001001;
  /* TG68KdotC_Kernel.vhd:3896:50  */
  assign n8912_o = opcode[6];
  assign n8914_o = n7915_o[1];
  assign n8915_o = n7897_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8916_o = n2184_o ? n8914_o : n8915_o;
  /* TG68KdotC_Kernel.vhd:3896:41  */
  assign n8917_o = n8912_o ? 1'b1 : n8916_o;
  /* TG68KdotC_Kernel.vhd:3899:50  */
  assign n8918_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3899:53  */
  assign n8919_o = ~n8918_o;
  /* TG68KdotC_Kernel.vhd:3899:41  */
  assign n8922_o = n8919_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3891:33  */
  assign n8924_o = micro_state == 7'b1001010;
  /* TG68KdotC_Kernel.vhd:3906:50  */
  assign n8925_o = opcode[6];
  assign n8928_o = n7915_o[3];
  assign n8929_o = n7897_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8930_o = n2184_o ? n8928_o : n8929_o;
  /* TG68KdotC_Kernel.vhd:3906:41  */
  assign n8931_o = n8925_o ? 1'b1 : n8930_o;
  assign n8932_o = n7919_o[9];
  assign n8933_o = n7899_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8934_o = n2184_o ? n8932_o : n8933_o;
  /* TG68KdotC_Kernel.vhd:3906:41  */
  assign n8935_o = n8925_o ? 1'b1 : n8934_o;
  /* TG68KdotC_Kernel.vhd:3910:50  */
  assign n8936_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3910:53  */
  assign n8937_o = ~n8936_o;
  /* TG68KdotC_Kernel.vhd:3910:41  */
  assign n8940_o = n8937_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3905:33  */
  assign n8942_o = micro_state == 7'b1001011;
  /* TG68KdotC_Kernel.vhd:3917:50  */
  assign n8943_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:3921:58  */
  assign n8947_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3921:61  */
  assign n8948_o = ~n8947_o;
  /* TG68KdotC_Kernel.vhd:3921:49  */
  assign n8951_o = n8948_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8953_o = n8943_o ? n7805_o : 2'b01;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8954_o = n8943_o ? n8951_o : n8058_o;
  assign n8955_o = n7915_o[3];
  assign n8956_o = n7897_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8957_o = n2184_o ? n8955_o : n8956_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8958_o = n8943_o ? 1'b1 : n8957_o;
  assign n8959_o = n7919_o[9];
  assign n8960_o = n7899_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8961_o = n2184_o ? n8959_o : n8960_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8962_o = n8943_o ? 1'b1 : n8961_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8963_o = n8943_o ? 1'b1 : n7951_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8965_o = n8943_o ? 7'b1001101 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3916:33  */
  assign n8967_o = micro_state == 7'b1001100;
  /* TG68KdotC_Kernel.vhd:3931:50  */
  assign n8968_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3931:53  */
  assign n8969_o = ~n8968_o;
  /* TG68KdotC_Kernel.vhd:3931:41  */
  assign n8972_o = n8969_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3930:33  */
  assign n8974_o = micro_state == 7'b1001101;
  /* TG68KdotC_Kernel.vhd:3937:33  */
  assign n8976_o = micro_state == 7'b1001110;
  /* TG68KdotC_Kernel.vhd:3941:50  */
  assign n8977_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3941:59  */
  assign n8979_o = n8977_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3941:41  */
  assign n8982_o = n8979_o ? 6'b001110 : 6'b011110;
  /* TG68KdotC_Kernel.vhd:3940:33  */
  assign n8984_o = micro_state == 7'b1010001;
  /* TG68KdotC_Kernel.vhd:3950:51  */
  assign n8987_o = rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:3950:41  */
  assign n8990_o = n8987_o ? 7'b1010011 : 7'b1010010;
  /* TG68KdotC_Kernel.vhd:3948:33  */
  assign n8992_o = micro_state == 7'b1010010;
  /* TG68KdotC_Kernel.vhd:3957:50  */
  assign n8993_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3957:54  */
  assign n8994_o = ~n8993_o;
  /* TG68KdotC_Kernel.vhd:3957:41  */
  assign n8996_o = n8994_o ? 1'b1 : n7934_o;
  /* TG68KdotC_Kernel.vhd:3962:50  */
  assign n8998_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3962:54  */
  assign n8999_o = ~n8998_o;
  /* TG68KdotC_Kernel.vhd:3962:59  */
  assign n9001_o = 1'b1 & n8999_o;
  /* TG68KdotC_Kernel.vhd:3965:58  */
  assign n9003_o = sndopc[10];
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n9005_o = n9009_o ? 2'b01 : n8058_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n9007_o = n9017_o ? 7'b1010100 : n8074_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n9009_o = n9003_o & n9001_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n9011_o = n9001_o ? 1'b1 : n7845_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n9012_o = n9001_o ? 1'b1 : n7913_o;
  assign n9013_o = n7922_o[4];
  assign n9014_o = n7715_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9015_o = n2184_o ? n9013_o : n9014_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n9016_o = n9001_o ? 1'b1 : n9015_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n9017_o = n9003_o & n9001_o;
  /* TG68KdotC_Kernel.vhd:3956:33  */
  assign n9019_o = micro_state == 7'b1010011;
  /* TG68KdotC_Kernel.vhd:3972:33  */
  assign n9024_o = micro_state == 7'b1010100;
  /* TG68KdotC_Kernel.vhd:3978:33  */
  assign n9026_o = micro_state == 7'b1010101;
  /* TG68KdotC_Kernel.vhd:3982:51  */
  assign n9027_o = op2out[31:16];
  /* TG68KdotC_Kernel.vhd:3982:65  */
  assign n9029_o = n9027_o == 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3982:83  */
  assign n9030_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3982:74  */
  assign n9031_o = n9029_o | n9030_o;
  /* TG68KdotC_Kernel.vhd:3982:92  */
  assign n9033_o = n9031_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3982:117  */
  assign n9034_o = op2out[15:0];
  /* TG68KdotC_Kernel.vhd:3982:130  */
  assign n9036_o = n9034_o == 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3982:107  */
  assign n9037_o = n9036_o & n9033_o;
  /* TG68KdotC_Kernel.vhd:3982:41  */
  assign n9040_o = n9037_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3982:41  */
  assign n9042_o = n9037_o ? n8074_o : 7'b1010111;
  /* TG68KdotC_Kernel.vhd:3981:33  */
  assign n9045_o = micro_state == 7'b1010110;
  /* TG68KdotC_Kernel.vhd:3990:50  */
  assign n9046_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3990:59  */
  assign n9048_o = n9046_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3990:41  */
  assign n9051_o = n9048_o ? 6'b001101 : 6'b011101;
  /* TG68KdotC_Kernel.vhd:3989:33  */
  assign n9053_o = micro_state == 7'b1010111;
  /* TG68KdotC_Kernel.vhd:3999:51  */
  assign n9056_o = rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:3999:41  */
  assign n9059_o = n9056_o ? 7'b1011001 : 7'b1011000;
  /* TG68KdotC_Kernel.vhd:3997:33  */
  assign n9061_o = micro_state == 7'b1011000;
  /* TG68KdotC_Kernel.vhd:4005:51  */
  assign n9062_o = ~z_error;
  /* TG68KdotC_Kernel.vhd:4005:70  */
  assign n9063_o = ~set_v_flag;
  /* TG68KdotC_Kernel.vhd:4005:56  */
  assign n9064_o = n9063_o & n9062_o;
  /* TG68KdotC_Kernel.vhd:4005:41  */
  assign n9066_o = n9064_o ? 1'b1 : n7913_o;
  /* TG68KdotC_Kernel.vhd:4008:50  */
  assign n9067_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:4008:54  */
  assign n9068_o = ~n9067_o;
  /* TG68KdotC_Kernel.vhd:4008:59  */
  assign n9070_o = 1'b1 & n9068_o;
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n9073_o = n9070_o ? 2'b01 : n8058_o;
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n9076_o = n9070_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n9077_o = n9070_o ? 1'b1 : n7950_o;
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n9079_o = n9070_o ? 7'b1011010 : n8074_o;
  /* TG68KdotC_Kernel.vhd:4004:33  */
  assign n9082_o = micro_state == 7'b1011001;
  /* TG68KdotC_Kernel.vhd:4017:48  */
  assign n9083_o = exec[34];
  /* TG68KdotC_Kernel.vhd:4017:41  */
  assign n9086_o = n9083_o ? 1'b1 : n7913_o;
  assign n9087_o = n7919_o[3];
  assign n9088_o = n7899_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9089_o = n2184_o ? n9087_o : n9088_o;
  /* TG68KdotC_Kernel.vhd:4017:41  */
  assign n9090_o = n9083_o ? n9089_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4016:33  */
  assign n9093_o = micro_state == 7'b1011010;
  /* TG68KdotC_Kernel.vhd:4026:50  */
  assign n9094_o = op2out[5:0];
  /* TG68KdotC_Kernel.vhd:4026:62  */
  assign n9096_o = n9094_o != 6'b000000;
  /* TG68KdotC_Kernel.vhd:4027:70  */
  assign n9097_o = op2out[5:0];
  /* TG68KdotC_Kernel.vhd:4026:41  */
  assign n9099_o = n9096_o ? n9097_o : n7851_o;
  assign n9100_o = n7982_o[23];
  /* TG68KdotC_Kernel.vhd:4026:41  */
  assign n9101_o = n9096_o ? n9100_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4025:33  */
  assign n9103_o = micro_state == 7'b1001111;
  /* TG68KdotC_Kernel.vhd:4032:33  */
  assign n9105_o = micro_state == 7'b1010000;
  assign n9106_o = {n9105_o, n9103_o, n9093_o, n9082_o, n9061_o, n9053_o, n9045_o, n9026_o, n9024_o, n9019_o, n8992_o, n8984_o, n8976_o, n8974_o, n8967_o, n8942_o, n8924_o, n8908_o, n8863_o, n8860_o, n8858_o, n8856_o, n8839_o, n8837_o, n8822_o, n8808_o, n8805_o, n8802_o, n8799_o, n8796_o, n8793_o, n8790_o, n8787_o, n8783_o, n8780_o, n8774_o, n8758_o, n8755_o, n8752_o, n8749_o, n8746_o, n8742_o, n8734_o, n8726_o, n8724_o, n8709_o, n8699_o, n8692_o, n8664_o, n8638_o, n8634_o, n8630_o, n8587_o, n8584_o, n8572_o, n8569_o, n8563_o, n8559_o, n8532_o, n8530_o, n8525_o, n8523_o, n8505_o, n8486_o, n8480_o, n8462_o, n8460_o, n8453_o, n8451_o, n8442_o, n8423_o, n8405_o, n8401_o, n8352_o, n8349_o, n8303_o, n8301_o, n8281_o, n8264_o, n8261_o, n8212_o, n8209_o, n8158_o, n8155_o, n8152_o};
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9109_o = 1'b1;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9109_o = n8466_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9109_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9109_o = n8444_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9109_o = n7804_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9109_o = n7804_o;
      default: n9109_o = n7804_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n8953_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9126_o = n8846_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b01;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b01;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9126_o = 2'b01;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9126_o = n8767_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9126_o = 2'b10;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9126_o = n8721_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9126_o = n7805_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9126_o = n7805_o;
      default: n9126_o = n7805_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9127_o = n8509_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9127_o = n8495_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9127_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9127_o = n7806_o;
      default: n9127_o = n7806_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n9073_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n9005_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8972_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8954_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8940_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8922_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9169_o = n8848_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9169_o = n8829_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9169_o = n8679_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9169_o = n8655_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9169_o = n8598_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9169_o = n8540_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9169_o = n8519_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9169_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9169_o = n8436_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9169_o = n8417_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9169_o = n8389_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9169_o = n8332_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9169_o = n8293_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9169_o = n8275_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9169_o = 2'b10;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9169_o = n8249_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9169_o = n8191_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9169_o = n8058_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9169_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9169_o = n8058_o;
      default: n9169_o = n8058_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9172_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9172_o = n8251_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9172_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9172_o = 1'b0;
      default: n9172_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9175_o = n8475_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9175_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9175_o = 1'b0;
      default: n9175_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9180_o = n8697_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9180_o = n8295_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9180_o = n8252_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9180_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9180_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9180_o = n7808_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9180_o = 1'b1;
      default: n9180_o = n7808_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9182_o = n8335_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9182_o = n8194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9182_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9182_o = 1'b0;
      default: n9182_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9192_o = n8428_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9192_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9192_o = n8356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9192_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9192_o = n8338_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9192_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9192_o = n8285_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9192_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9192_o = n8216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9192_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9192_o = n8197_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9192_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9192_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9192_o = 1'b0;
      default: n9192_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9196_o = n8477_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9196_o = n8457_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9196_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9196_o = n8447_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9196_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9196_o = 1'b0;
      default: n9196_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9214_o = n8850_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9214_o = n8831_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9214_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9214_o = n7819_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9214_o = n7819_o;
      default: n9214_o = n7819_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9216_o = n8777_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9216_o = n8768_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9216_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9216_o = n8137_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9216_o = n8137_o;
      default: n9216_o = n8137_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b1;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9219_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9219_o = 1'b0;
      default: n9219_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9222_o = 1'b1;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9222_o = n8031_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9222_o = n8031_o;
      default: n9222_o = n8031_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9225_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9225_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9225_o = 1'b0;
      default: n9225_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9229_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9229_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9229_o = 1'b0;
      default: n9229_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9233_o = n8601_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9233_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9233_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9233_o = 1'b0;
      default: n9233_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9236_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9236_o = n7839_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9236_o = n7839_o;
      default: n9236_o = n7839_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9241_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9241_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9241_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9241_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9241_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9241_o = n8060_o;
      default: n9241_o = n8060_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9243_o = n8603_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9243_o = n8560_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9243_o = n8512_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9243_o = n8498_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9243_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9243_o = 1'b0;
      default: n9243_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9248_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9248_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9248_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9248_o = 1'b0;
      default: n9248_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9251_o = n8606_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9251_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9251_o = 1'b0;
      default: n9251_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = 1'b1;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n9011_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9257_o = n8608_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9257_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9257_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9257_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9257_o = n7845_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9257_o = n7845_o;
      default: n9257_o = n7845_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = n9076_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9261_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9261_o = n8543_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9261_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9261_o = 1'b0;
      default: n9261_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9266_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9266_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9266_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9266_o = n8100_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9266_o = n8100_o;
      default: n9266_o = n8100_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n9099_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n9051_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n8982_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9267_o = n7851_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9267_o = n7851_o;
      default: n9267_o = n7851_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9271_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9271_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9271_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9271_o = n7855_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9271_o = n7855_o;
      default: n9271_o = n7855_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9274_o = 1'b1;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9274_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9274_o = 1'b0;
      default: n9274_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9278_o = 1'b1;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9278_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9278_o = 1'b0;
      default: n9278_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n8903_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9280_o = n7857_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9280_o = n7857_o;
      default: n9280_o = n7857_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8905_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9281_o = n8528_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9281_o = n8140_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9281_o = n8140_o;
      default: n9281_o = n8140_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9284_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9284_o = n8339_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9284_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9284_o = n8198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9284_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9284_o = n2157_o;
      default: n9284_o = n2157_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = n9040_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9286_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9286_o = 1'b0;
      default: n9286_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9288_o = 1'b1;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9288_o = n7903_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9288_o = n7903_o;
      default: n9288_o = n7903_o;
    endcase
  assign n9289_o = n1909_o[20];
  assign n9290_o = n7896_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9291_o = n2184_o ? n9289_o : n9290_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = 1'b1;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9292_o = n9291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9292_o = n9291_o;
      default: n9292_o = n9291_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = 1'b1;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = 1'b1;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9293_o = n7938_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9293_o = n7938_o;
      default: n9293_o = n7938_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9294_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9294_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9294_o = n8199_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9294_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9294_o = n2164_o;
      default: n9294_o = n2164_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = 1'b1;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9295_o = n7907_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9295_o = n7907_o;
      default: n9295_o = n7907_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9296_o = n8769_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9296_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9296_o = n1960_o;
      default: n9296_o = n1960_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9297_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9297_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9297_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9297_o = n7909_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9297_o = n7909_o;
      default: n9297_o = n7909_o;
    endcase
  assign n9298_o = n1909_o[27];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9299_o = 1'b1;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9299_o = 1'b1;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9299_o = n8610_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9299_o = n8545_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9299_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9299_o = n9298_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9299_o = n9298_o;
      default: n9299_o = n9298_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n9086_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n9066_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n9012_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9300_o = n8901_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9300_o = 1'b1;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9300_o = 1'b1;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9300_o = n8648_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9300_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9300_o = n8611_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9300_o = n8546_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9300_o = n7913_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9300_o = n7913_o;
      default: n9300_o = n7913_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9301_o = 1'b1;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9301_o = n8816_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9301_o = n7946_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9301_o = n7946_o;
      default: n9301_o = n7946_o;
    endcase
  assign n9302_o = n7915_o[1];
  assign n9303_o = n7897_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9304_o = n2184_o ? n9302_o : n9303_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n8917_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9305_o = n9304_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9305_o = n9304_o;
      default: n9305_o = n9304_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9306_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9306_o = n8104_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9306_o = n8104_o;
      default: n9306_o = n8104_o;
    endcase
  assign n9307_o = n7915_o[3];
  assign n9308_o = n7897_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9309_o = n2184_o ? n9307_o : n9308_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n8958_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n8931_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9310_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9310_o = n9309_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9310_o = n9309_o;
      default: n9310_o = n9309_o;
    endcase
  assign n9311_o = n7915_o[4];
  assign n9312_o = n7897_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9313_o = n2184_o ? n9311_o : n9312_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9314_o = n8683_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9314_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9314_o = n8615_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9314_o = n8550_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9314_o = n9313_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9314_o = n9313_o;
      default: n9314_o = n9313_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9315_o = n7947_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9315_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9315_o = 1'b1;
      default: n9315_o = n7947_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9316_o = n8851_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9316_o = n8832_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9316_o = 1'b1;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9316_o = 1'b1;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9316_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9316_o = n8124_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9316_o = n8124_o;
      default: n9316_o = n8124_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9317_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9317_o = n8108_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9317_o = n8108_o;
      default: n9317_o = n8108_o;
    endcase
  assign n9318_o = n7919_o[3];
  assign n9319_o = n7899_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9320_o = n2184_o ? n9318_o : n9319_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9090_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9321_o = n9320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9321_o = n9320_o;
      default: n9321_o = n9320_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9322_o = n8739_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9322_o = n8731_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9322_o = n8714_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9322_o = n8704_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9322_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9322_o = n8112_o;
      default: n9322_o = n8112_o;
    endcase
  assign n9323_o = n7919_o[9];
  assign n9324_o = n7899_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9325_o = n2184_o ? n9323_o : n9324_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n8962_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n8935_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9326_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9326_o = n8687_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9326_o = n8660_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9326_o = n9325_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9326_o = n9325_o;
      default: n9326_o = n9325_o;
    endcase
  assign n9327_o = n7919_o[10];
  assign n9328_o = n7899_o[10];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9329_o = n2184_o ? n9327_o : n9328_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9330_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9330_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9330_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9330_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9330_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9330_o = n9329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9330_o = n9329_o;
      default: n9330_o = n9329_o;
    endcase
  assign n9331_o = n7919_o[11];
  assign n9332_o = n7899_o[11];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9333_o = n2184_o ? n9331_o : n9332_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9334_o = 1'b1;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9334_o = 1'b1;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9334_o = n9333_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9334_o = n9333_o;
      default: n9334_o = n9333_o;
    endcase
  assign n9335_o = n7919_o[12];
  assign n9336_o = n7899_o[12];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9337_o = n2184_o ? n9335_o : n9336_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9338_o = n8820_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9338_o = 1'b1;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9338_o = n9337_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9338_o = n9337_o;
      default: n9338_o = n9337_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9339_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9339_o = n8616_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9339_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9339_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9339_o = n8296_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9339_o = n8253_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9339_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9339_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9339_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9339_o = 1'b1;
      default: n9339_o = n2170_o;
    endcase
  assign n9340_o = n7922_o[1];
  assign n9341_o = n7715_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9342_o = n2184_o ? n9340_o : n9341_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9343_o = n8620_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9343_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9343_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9343_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9343_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9343_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9343_o = n8393_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9343_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9343_o = n9342_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9343_o = n9342_o;
      default: n9343_o = n9342_o;
    endcase
  assign n9344_o = n7922_o[4];
  assign n9345_o = n7715_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9346_o = n2184_o ? n9344_o : n9345_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9016_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9347_o = n9346_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9347_o = n9346_o;
      default: n9347_o = n9346_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n9077_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9348_o = n7950_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9348_o = n7950_o;
      default: n9348_o = n7950_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9349_o = n8688_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9349_o = n7925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9349_o = n7925_o;
      default: n9349_o = n7925_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9350_o = 1'b1;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9350_o = n8437_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9350_o = n8394_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9350_o = n8340_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9350_o = n8297_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9350_o = n8254_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9350_o = n8200_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9350_o = n7952_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9350_o = n7952_o;
      default: n9350_o = n7952_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n8963_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9351_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9351_o = n7951_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9351_o = n7951_o;
      default: n9351_o = n7951_o;
    endcase
  assign n9352_o = n7929_o[0];
  assign n9353_o = n7900_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9354_o = n2184_o ? n9352_o : n9353_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9355_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9355_o = n8421_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9355_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9355_o = n8398_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9355_o = n8344_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9355_o = n8279_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9355_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9355_o = n8258_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9355_o = n8204_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9355_o = n9354_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9355_o = n9354_o;
      default: n9355_o = n9354_o;
    endcase
  assign n9356_o = n1909_o[79];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9357_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9357_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9357_o = n9356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9357_o = n9356_o;
      default: n9357_o = n9356_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n8996_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9358_o = n8621_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9358_o = n7934_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9358_o = n7934_o;
      default: n9358_o = n7934_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9359_o = n8551_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9359_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9359_o = n1925_o;
      default: n9359_o = n1925_o;
    endcase
  assign n9360_o = n1909_o[84];
  assign n9361_o = n7901_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9362_o = n2184_o ? n9360_o : n9361_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9363_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9363_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9363_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9363_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9363_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9363_o = n9362_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9363_o = n9362_o;
      default: n9363_o = n9362_o;
    endcase
  assign n9364_o = n1909_o[85];
  assign n9365_o = n7901_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9366_o = n2184_o ? n9364_o : n9365_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9367_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9367_o = n8625_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9367_o = n8555_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9367_o = n9366_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9367_o = n9366_o;
      default: n9367_o = n9366_o;
    endcase
  assign n9368_o = n1909_o[86];
  assign n9369_o = n7901_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9370_o = n2184_o ? n9368_o : n9369_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9371_o = n8578_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9371_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9371_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9371_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9371_o = n9370_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9371_o = n9370_o;
      default: n9371_o = n9370_o;
    endcase
  assign n9372_o = n1909_o[87];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9373_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9373_o = n9372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9373_o = n9372_o;
      default: n9373_o = n9372_o;
    endcase
  assign n9374_o = n1909_o[88];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9375_o = n8516_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9375_o = n8493_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9375_o = n9374_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9375_o = n9374_o;
      default: n9375_o = n9374_o;
    endcase
  assign n9376_o = n1909_o[19:17];
  assign n9377_o = n7896_o[2:0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9378_o = n2184_o ? n9376_o : n9377_o;
  assign n9379_o = n1909_o[28];
  assign n9380_o = n7915_o[0];
  assign n9381_o = n7897_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9382_o = n2184_o ? n9380_o : n9381_o;
  assign n9386_o = n7919_o[2];
  assign n9387_o = n7899_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9388_o = n2184_o ? n9386_o : n9387_o;
  assign n9392_o = n7919_o[8:5];
  assign n9393_o = n7899_o[8:5];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9394_o = n2184_o ? n9392_o : n9393_o;
  assign n9401_o = n7919_o[15:13];
  assign n9402_o = n7899_o[15:13];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9403_o = n2184_o ? n9401_o : n9402_o;
  assign n9407_o = n7922_o[0];
  assign n9408_o = n7715_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9409_o = n2184_o ? n9407_o : n9408_o;
  assign n9410_o = n7922_o[3:2];
  assign n9411_o = n7715_o[3:2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9412_o = n2184_o ? n9410_o : n9411_o;
  assign n9413_o = n7929_o[1];
  assign n9414_o = n7900_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9415_o = n2184_o ? n9413_o : n9414_o;
  assign n9416_o = n1909_o[78:75];
  assign n9424_o = n7982_o[23];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9101_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9425_o = n9424_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9425_o = n9424_o;
      default: n9425_o = n9424_o;
    endcase
  assign n9426_o = n7982_o[25:24];
  assign n9427_o = n7982_o[22:21];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n9106_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n9079_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n9059_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1011000;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n9042_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1010110;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n9007_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8990_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1010010;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1001110;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8965_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1001100;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1001011;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b0110001;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b0000001;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9473_o = n8854_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b0101110;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9473_o = n8835_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b0101100;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b0110011;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1011110;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1011101;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1011100;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1011011;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9473_o = 7'b1001000;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9473_o = 7'b1000111;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9473_o = 7'b0011000;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9473_o = 7'b0110110;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9473_o = 7'b0110101;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9473_o = n8772_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9473_o = 7'b0110011;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9473_o = 7'b0100110;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9473_o = 7'b0100100;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9473_o = 7'b0100000;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9473_o = 7'b0011111;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9473_o = n8690_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9473_o = n8662_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9473_o = 7'b0011000;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9473_o = n8628_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9473_o = 7'b0111110;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9473_o = 7'b0111101;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9473_o = 7'b0111100;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9473_o = 7'b0111011;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9473_o = 7'b0111010;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9473_o = n8557_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9473_o = 7'b0111000;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9473_o = 7'b1000101;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9473_o = n8521_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9473_o = 7'b1000011;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9473_o = 7'b1000010;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9473_o = n8471_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9473_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9473_o = 7'b0011000;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9473_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9473_o = n8449_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9473_o = n8440_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9473_o = 7'b0010010;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9473_o = 7'b0010001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9473_o = n8399_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9473_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9473_o = n8347_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9473_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9473_o = n8299_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9473_o = 7'b0001110;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9473_o = 7'b0001101;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9473_o = n8259_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9473_o = n8207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9473_o = n8074_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9473_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9473_o = n8074_o;
      default: n9473_o = n8074_o;
    endcase
  /* TG68KdotC_Kernel.vhd:4049:41  */
  assign n9478_o = exec[33];
  /* TG68KdotC_Kernel.vhd:4049:33  */
  assign n9479_o = n9478_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:4050:27  */
  assign n9480_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:4051:47  */
  assign n9481_o = reg_qa[2:0];
  /* TG68KdotC_Kernel.vhd:4051:19  */
  assign n9483_o = n9480_o == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:4052:47  */
  assign n9484_o = reg_qa[2:0];
  /* TG68KdotC_Kernel.vhd:4052:19  */
  assign n9486_o = n9480_o == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:4053:48  */
  assign n9487_o = reg_qa[3:0];
  /* TG68KdotC_Kernel.vhd:4053:19  */
  assign n9489_o = n9480_o == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:4054:19  */
  assign n9491_o = n9480_o == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:4055:19  */
  assign n9493_o = n9480_o == 12'b100000000001;
  /* TG68KdotC_Kernel.vhd:4056:19  */
  assign n9495_o = n9480_o == 12'b100000000010;
  /* TG68KdotC_Kernel.vhd:4057:19  */
  assign n9497_o = n9480_o == 12'b100000000011;
  /* TG68KdotC_Kernel.vhd:4058:19  */
  assign n9499_o = n9480_o == 12'b100000000100;
  assign n9500_o = {n9499_o, n9497_o, n9495_o, n9493_o, n9491_o, n9489_o, n9486_o, n9483_o};
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9500_o)
      8'b10000000: n9501_o = vbr;
      8'b01000000: n9501_o = vbr;
      8'b00100000: n9501_o = vbr;
      8'b00010000: n9501_o = reg_qa;
      8'b00001000: n9501_o = vbr;
      8'b00000100: n9501_o = vbr;
      8'b00000010: n9501_o = vbr;
      8'b00000001: n9501_o = vbr;
      default: n9501_o = vbr;
    endcase
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9500_o)
      8'b10000000: n9502_o = cacr;
      8'b01000000: n9502_o = cacr;
      8'b00100000: n9502_o = cacr;
      8'b00010000: n9502_o = cacr;
      8'b00001000: n9502_o = cacr;
      8'b00000100: n9502_o = n9487_o;
      8'b00000010: n9502_o = cacr;
      8'b00000001: n9502_o = cacr;
      default: n9502_o = cacr;
    endcase
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9500_o)
      8'b10000000: n9503_o = dfc;
      8'b01000000: n9503_o = dfc;
      8'b00100000: n9503_o = dfc;
      8'b00010000: n9503_o = dfc;
      8'b00001000: n9503_o = dfc;
      8'b00000100: n9503_o = dfc;
      8'b00000010: n9503_o = n9484_o;
      8'b00000001: n9503_o = dfc;
      default: n9503_o = dfc;
    endcase
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9500_o)
      8'b10000000: n9504_o = sfc;
      8'b01000000: n9504_o = sfc;
      8'b00100000: n9504_o = sfc;
      8'b00010000: n9504_o = sfc;
      8'b00001000: n9504_o = sfc;
      8'b00000100: n9504_o = sfc;
      8'b00000010: n9504_o = sfc;
      8'b00000001: n9504_o = n9481_o;
      default: n9504_o = sfc;
    endcase
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9505_o = n9479_o ? n9501_o : vbr;
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9506_o = n9479_o ? n9502_o : cacr;
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9507_o = n9479_o ? n9503_o : dfc;
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9508_o = n9479_o ? n9504_o : sfc;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9510_o = reset ? 32'b00000000000000000000000000000000 : n9505_o;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9512_o = reset ? 4'b0000 : n9506_o;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9513_o = reset ? dfc : n9507_o;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9514_o = reset ? sfc : n9508_o;
  /* TG68KdotC_Kernel.vhd:4065:19  */
  assign n9519_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:4066:78  */
  assign n9521_o = {29'b00000000000000000000000000000, sfc};
  /* TG68KdotC_Kernel.vhd:4066:17  */
  assign n9523_o = n9519_o == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:4067:78  */
  assign n9525_o = {29'b00000000000000000000000000000, dfc};
  /* TG68KdotC_Kernel.vhd:4067:17  */
  assign n9527_o = n9519_o == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:4068:79  */
  assign n9529_o = cacr & 4'b0011;
  /* TG68KdotC_Kernel.vhd:4068:71  */
  assign n9531_o = {28'b0000000000000000000000000000, n9529_o};
  /* TG68KdotC_Kernel.vhd:4068:11  */
  assign n9533_o = n9519_o == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:4070:11  */
  assign n9535_o = n9519_o == 12'b100000000001;
  assign n9536_o = {n9535_o, n9533_o, n9527_o, n9523_o};
  /* TG68KdotC_Kernel.vhd:4065:9  */
  always @*
    case (n9536_o)
      4'b1000: n9538_o = vbr;
      4'b0100: n9538_o = n9531_o;
      4'b0010: n9538_o = n9525_o;
      4'b0001: n9538_o = n9521_o;
      default: n9538_o = 32'b00000000000000000000000000000000;
    endcase
  /* TG68KdotC_Kernel.vhd:4084:32  */
  assign n9543_o = exe_opcode[11:8];
  /* TG68KdotC_Kernel.vhd:4085:25  */
  assign n9545_o = n9543_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4086:25  */
  assign n9547_o = n9543_o == 4'b0001;
  /* TG68KdotC_Kernel.vhd:4087:65  */
  assign n9548_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4087:56  */
  assign n9549_o = ~n9548_o;
  /* TG68KdotC_Kernel.vhd:4087:82  */
  assign n9550_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4087:73  */
  assign n9551_o = ~n9550_o;
  /* TG68KdotC_Kernel.vhd:4087:69  */
  assign n9552_o = n9549_o & n9551_o;
  /* TG68KdotC_Kernel.vhd:4087:25  */
  assign n9554_o = n9543_o == 4'b0010;
  /* TG68KdotC_Kernel.vhd:4088:60  */
  assign n9555_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4088:72  */
  assign n9556_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4088:64  */
  assign n9557_o = n9555_o | n9556_o;
  /* TG68KdotC_Kernel.vhd:4088:25  */
  assign n9559_o = n9543_o == 4'b0011;
  /* TG68KdotC_Kernel.vhd:4089:64  */
  assign n9560_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4089:55  */
  assign n9561_o = ~n9560_o;
  /* TG68KdotC_Kernel.vhd:4089:25  */
  assign n9563_o = n9543_o == 4'b0100;
  /* TG68KdotC_Kernel.vhd:4090:60  */
  assign n9564_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4090:25  */
  assign n9566_o = n9543_o == 4'b0101;
  /* TG68KdotC_Kernel.vhd:4091:64  */
  assign n9567_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4091:55  */
  assign n9568_o = ~n9567_o;
  /* TG68KdotC_Kernel.vhd:4091:25  */
  assign n9570_o = n9543_o == 4'b0110;
  /* TG68KdotC_Kernel.vhd:4092:60  */
  assign n9571_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4092:25  */
  assign n9573_o = n9543_o == 4'b0111;
  /* TG68KdotC_Kernel.vhd:4093:64  */
  assign n9574_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4093:55  */
  assign n9575_o = ~n9574_o;
  /* TG68KdotC_Kernel.vhd:4093:25  */
  assign n9577_o = n9543_o == 4'b1000;
  /* TG68KdotC_Kernel.vhd:4094:60  */
  assign n9578_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4094:25  */
  assign n9580_o = n9543_o == 4'b1001;
  /* TG68KdotC_Kernel.vhd:4095:64  */
  assign n9581_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4095:55  */
  assign n9582_o = ~n9581_o;
  /* TG68KdotC_Kernel.vhd:4095:25  */
  assign n9584_o = n9543_o == 4'b1010;
  /* TG68KdotC_Kernel.vhd:4096:60  */
  assign n9585_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4096:25  */
  assign n9587_o = n9543_o == 4'b1011;
  /* TG68KdotC_Kernel.vhd:4097:61  */
  assign n9588_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4097:74  */
  assign n9589_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4097:65  */
  assign n9590_o = n9588_o & n9589_o;
  /* TG68KdotC_Kernel.vhd:4097:92  */
  assign n9591_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4097:83  */
  assign n9592_o = ~n9591_o;
  /* TG68KdotC_Kernel.vhd:4097:109  */
  assign n9593_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4097:100  */
  assign n9594_o = ~n9593_o;
  /* TG68KdotC_Kernel.vhd:4097:96  */
  assign n9595_o = n9592_o & n9594_o;
  /* TG68KdotC_Kernel.vhd:4097:79  */
  assign n9596_o = n9590_o | n9595_o;
  /* TG68KdotC_Kernel.vhd:4097:25  */
  assign n9598_o = n9543_o == 4'b1100;
  /* TG68KdotC_Kernel.vhd:4098:61  */
  assign n9599_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4098:78  */
  assign n9600_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4098:69  */
  assign n9601_o = ~n9600_o;
  /* TG68KdotC_Kernel.vhd:4098:65  */
  assign n9602_o = n9599_o & n9601_o;
  /* TG68KdotC_Kernel.vhd:4098:96  */
  assign n9603_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4098:87  */
  assign n9604_o = ~n9603_o;
  /* TG68KdotC_Kernel.vhd:4098:109  */
  assign n9605_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4098:100  */
  assign n9606_o = n9604_o & n9605_o;
  /* TG68KdotC_Kernel.vhd:4098:83  */
  assign n9607_o = n9602_o | n9606_o;
  /* TG68KdotC_Kernel.vhd:4098:25  */
  assign n9609_o = n9543_o == 4'b1101;
  /* TG68KdotC_Kernel.vhd:4099:61  */
  assign n9610_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4099:74  */
  assign n9611_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4099:65  */
  assign n9612_o = n9610_o & n9611_o;
  /* TG68KdotC_Kernel.vhd:4099:91  */
  assign n9613_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4099:82  */
  assign n9614_o = ~n9613_o;
  /* TG68KdotC_Kernel.vhd:4099:78  */
  assign n9615_o = n9612_o & n9614_o;
  /* TG68KdotC_Kernel.vhd:4099:109  */
  assign n9616_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4099:100  */
  assign n9617_o = ~n9616_o;
  /* TG68KdotC_Kernel.vhd:4099:126  */
  assign n9618_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4099:117  */
  assign n9619_o = ~n9618_o;
  /* TG68KdotC_Kernel.vhd:4099:113  */
  assign n9620_o = n9617_o & n9619_o;
  /* TG68KdotC_Kernel.vhd:4099:143  */
  assign n9621_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4099:134  */
  assign n9622_o = ~n9621_o;
  /* TG68KdotC_Kernel.vhd:4099:130  */
  assign n9623_o = n9620_o & n9622_o;
  /* TG68KdotC_Kernel.vhd:4099:96  */
  assign n9624_o = n9615_o | n9623_o;
  /* TG68KdotC_Kernel.vhd:4099:25  */
  assign n9626_o = n9543_o == 4'b1110;
  /* TG68KdotC_Kernel.vhd:4100:61  */
  assign n9627_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4100:78  */
  assign n9628_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4100:69  */
  assign n9629_o = ~n9628_o;
  /* TG68KdotC_Kernel.vhd:4100:65  */
  assign n9630_o = n9627_o & n9629_o;
  /* TG68KdotC_Kernel.vhd:4100:96  */
  assign n9631_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4100:87  */
  assign n9632_o = ~n9631_o;
  /* TG68KdotC_Kernel.vhd:4100:109  */
  assign n9633_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4100:100  */
  assign n9634_o = n9632_o & n9633_o;
  /* TG68KdotC_Kernel.vhd:4100:83  */
  assign n9635_o = n9630_o | n9634_o;
  /* TG68KdotC_Kernel.vhd:4100:122  */
  assign n9636_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4100:114  */
  assign n9637_o = n9635_o | n9636_o;
  /* TG68KdotC_Kernel.vhd:4100:25  */
  assign n9639_o = n9543_o == 4'b1111;
  assign n9640_o = {n9639_o, n9626_o, n9609_o, n9598_o, n9587_o, n9584_o, n9580_o, n9577_o, n9573_o, n9570_o, n9566_o, n9563_o, n9559_o, n9554_o, n9547_o, n9545_o};
  /* TG68KdotC_Kernel.vhd:4084:17  */
  always @*
    case (n9640_o)
      16'b1000000000000000: n9643_o = n9637_o;
      16'b0100000000000000: n9643_o = n9624_o;
      16'b0010000000000000: n9643_o = n9607_o;
      16'b0001000000000000: n9643_o = n9596_o;
      16'b0000100000000000: n9643_o = n9585_o;
      16'b0000010000000000: n9643_o = n9582_o;
      16'b0000001000000000: n9643_o = n9578_o;
      16'b0000000100000000: n9643_o = n9575_o;
      16'b0000000010000000: n9643_o = n9571_o;
      16'b0000000001000000: n9643_o = n9568_o;
      16'b0000000000100000: n9643_o = n9564_o;
      16'b0000000000010000: n9643_o = n9561_o;
      16'b0000000000001000: n9643_o = n9557_o;
      16'b0000000000000100: n9643_o = n9552_o;
      16'b0000000000000010: n9643_o = 1'b0;
      16'b0000000000000001: n9643_o = 1'b1;
      default: n9643_o = exe_condition;
    endcase
  /* TG68KdotC_Kernel.vhd:4112:54  */
  assign n9648_o = exec[69];
  /* TG68KdotC_Kernel.vhd:4114:60  */
  assign n9649_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:4115:43  */
  assign n9650_o = exec[69];
  /* TG68KdotC_Kernel.vhd:4115:68  */
  assign n9651_o = set[69];
  /* TG68KdotC_Kernel.vhd:4115:62  */
  assign n9652_o = n9650_o | n9651_o;
  /* TG68KdotC_Kernel.vhd:4117:49  */
  assign n9655_o = movem_regaddr == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4118:49  */
  assign n9658_o = movem_regaddr == 4'b0001;
  /* TG68KdotC_Kernel.vhd:4119:49  */
  assign n9661_o = movem_regaddr == 4'b0010;
  /* TG68KdotC_Kernel.vhd:4120:49  */
  assign n9664_o = movem_regaddr == 4'b0011;
  /* TG68KdotC_Kernel.vhd:4121:49  */
  assign n9667_o = movem_regaddr == 4'b0100;
  /* TG68KdotC_Kernel.vhd:4122:49  */
  assign n9670_o = movem_regaddr == 4'b0101;
  /* TG68KdotC_Kernel.vhd:4123:49  */
  assign n9673_o = movem_regaddr == 4'b0110;
  /* TG68KdotC_Kernel.vhd:4124:49  */
  assign n9676_o = movem_regaddr == 4'b0111;
  /* TG68KdotC_Kernel.vhd:4125:49  */
  assign n9679_o = movem_regaddr == 4'b1000;
  /* TG68KdotC_Kernel.vhd:4126:49  */
  assign n9682_o = movem_regaddr == 4'b1001;
  /* TG68KdotC_Kernel.vhd:4127:49  */
  assign n9685_o = movem_regaddr == 4'b1010;
  /* TG68KdotC_Kernel.vhd:4128:49  */
  assign n9688_o = movem_regaddr == 4'b1011;
  /* TG68KdotC_Kernel.vhd:4129:49  */
  assign n9691_o = movem_regaddr == 4'b1100;
  /* TG68KdotC_Kernel.vhd:4130:49  */
  assign n9694_o = movem_regaddr == 4'b1101;
  /* TG68KdotC_Kernel.vhd:4131:49  */
  assign n9697_o = movem_regaddr == 4'b1110;
  /* TG68KdotC_Kernel.vhd:4132:49  */
  assign n9700_o = movem_regaddr == 4'b1111;
  assign n9701_o = {n9700_o, n9697_o, n9694_o, n9691_o, n9688_o, n9685_o, n9682_o, n9679_o, n9676_o, n9673_o, n9670_o, n9667_o, n9664_o, n9661_o, n9658_o, n9655_o};
  assign n9702_o = sndopc[0];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9703_o = n9702_o;
      16'b0100000000000000: n9703_o = n9702_o;
      16'b0010000000000000: n9703_o = n9702_o;
      16'b0001000000000000: n9703_o = n9702_o;
      16'b0000100000000000: n9703_o = n9702_o;
      16'b0000010000000000: n9703_o = n9702_o;
      16'b0000001000000000: n9703_o = n9702_o;
      16'b0000000100000000: n9703_o = n9702_o;
      16'b0000000010000000: n9703_o = n9702_o;
      16'b0000000001000000: n9703_o = n9702_o;
      16'b0000000000100000: n9703_o = n9702_o;
      16'b0000000000010000: n9703_o = n9702_o;
      16'b0000000000001000: n9703_o = n9702_o;
      16'b0000000000000100: n9703_o = n9702_o;
      16'b0000000000000010: n9703_o = n9702_o;
      16'b0000000000000001: n9703_o = 1'b0;
      default: n9703_o = n9702_o;
    endcase
  assign n9704_o = sndopc[1];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9705_o = n9704_o;
      16'b0100000000000000: n9705_o = n9704_o;
      16'b0010000000000000: n9705_o = n9704_o;
      16'b0001000000000000: n9705_o = n9704_o;
      16'b0000100000000000: n9705_o = n9704_o;
      16'b0000010000000000: n9705_o = n9704_o;
      16'b0000001000000000: n9705_o = n9704_o;
      16'b0000000100000000: n9705_o = n9704_o;
      16'b0000000010000000: n9705_o = n9704_o;
      16'b0000000001000000: n9705_o = n9704_o;
      16'b0000000000100000: n9705_o = n9704_o;
      16'b0000000000010000: n9705_o = n9704_o;
      16'b0000000000001000: n9705_o = n9704_o;
      16'b0000000000000100: n9705_o = n9704_o;
      16'b0000000000000010: n9705_o = 1'b0;
      16'b0000000000000001: n9705_o = n9704_o;
      default: n9705_o = n9704_o;
    endcase
  assign n9706_o = sndopc[2];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9707_o = n9706_o;
      16'b0100000000000000: n9707_o = n9706_o;
      16'b0010000000000000: n9707_o = n9706_o;
      16'b0001000000000000: n9707_o = n9706_o;
      16'b0000100000000000: n9707_o = n9706_o;
      16'b0000010000000000: n9707_o = n9706_o;
      16'b0000001000000000: n9707_o = n9706_o;
      16'b0000000100000000: n9707_o = n9706_o;
      16'b0000000010000000: n9707_o = n9706_o;
      16'b0000000001000000: n9707_o = n9706_o;
      16'b0000000000100000: n9707_o = n9706_o;
      16'b0000000000010000: n9707_o = n9706_o;
      16'b0000000000001000: n9707_o = n9706_o;
      16'b0000000000000100: n9707_o = 1'b0;
      16'b0000000000000010: n9707_o = n9706_o;
      16'b0000000000000001: n9707_o = n9706_o;
      default: n9707_o = n9706_o;
    endcase
  assign n9708_o = sndopc[3];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9709_o = n9708_o;
      16'b0100000000000000: n9709_o = n9708_o;
      16'b0010000000000000: n9709_o = n9708_o;
      16'b0001000000000000: n9709_o = n9708_o;
      16'b0000100000000000: n9709_o = n9708_o;
      16'b0000010000000000: n9709_o = n9708_o;
      16'b0000001000000000: n9709_o = n9708_o;
      16'b0000000100000000: n9709_o = n9708_o;
      16'b0000000010000000: n9709_o = n9708_o;
      16'b0000000001000000: n9709_o = n9708_o;
      16'b0000000000100000: n9709_o = n9708_o;
      16'b0000000000010000: n9709_o = n9708_o;
      16'b0000000000001000: n9709_o = 1'b0;
      16'b0000000000000100: n9709_o = n9708_o;
      16'b0000000000000010: n9709_o = n9708_o;
      16'b0000000000000001: n9709_o = n9708_o;
      default: n9709_o = n9708_o;
    endcase
  assign n9710_o = sndopc[4];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9711_o = n9710_o;
      16'b0100000000000000: n9711_o = n9710_o;
      16'b0010000000000000: n9711_o = n9710_o;
      16'b0001000000000000: n9711_o = n9710_o;
      16'b0000100000000000: n9711_o = n9710_o;
      16'b0000010000000000: n9711_o = n9710_o;
      16'b0000001000000000: n9711_o = n9710_o;
      16'b0000000100000000: n9711_o = n9710_o;
      16'b0000000010000000: n9711_o = n9710_o;
      16'b0000000001000000: n9711_o = n9710_o;
      16'b0000000000100000: n9711_o = n9710_o;
      16'b0000000000010000: n9711_o = 1'b0;
      16'b0000000000001000: n9711_o = n9710_o;
      16'b0000000000000100: n9711_o = n9710_o;
      16'b0000000000000010: n9711_o = n9710_o;
      16'b0000000000000001: n9711_o = n9710_o;
      default: n9711_o = n9710_o;
    endcase
  assign n9712_o = sndopc[5];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9713_o = n9712_o;
      16'b0100000000000000: n9713_o = n9712_o;
      16'b0010000000000000: n9713_o = n9712_o;
      16'b0001000000000000: n9713_o = n9712_o;
      16'b0000100000000000: n9713_o = n9712_o;
      16'b0000010000000000: n9713_o = n9712_o;
      16'b0000001000000000: n9713_o = n9712_o;
      16'b0000000100000000: n9713_o = n9712_o;
      16'b0000000010000000: n9713_o = n9712_o;
      16'b0000000001000000: n9713_o = n9712_o;
      16'b0000000000100000: n9713_o = 1'b0;
      16'b0000000000010000: n9713_o = n9712_o;
      16'b0000000000001000: n9713_o = n9712_o;
      16'b0000000000000100: n9713_o = n9712_o;
      16'b0000000000000010: n9713_o = n9712_o;
      16'b0000000000000001: n9713_o = n9712_o;
      default: n9713_o = n9712_o;
    endcase
  assign n9714_o = sndopc[6];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9715_o = n9714_o;
      16'b0100000000000000: n9715_o = n9714_o;
      16'b0010000000000000: n9715_o = n9714_o;
      16'b0001000000000000: n9715_o = n9714_o;
      16'b0000100000000000: n9715_o = n9714_o;
      16'b0000010000000000: n9715_o = n9714_o;
      16'b0000001000000000: n9715_o = n9714_o;
      16'b0000000100000000: n9715_o = n9714_o;
      16'b0000000010000000: n9715_o = n9714_o;
      16'b0000000001000000: n9715_o = 1'b0;
      16'b0000000000100000: n9715_o = n9714_o;
      16'b0000000000010000: n9715_o = n9714_o;
      16'b0000000000001000: n9715_o = n9714_o;
      16'b0000000000000100: n9715_o = n9714_o;
      16'b0000000000000010: n9715_o = n9714_o;
      16'b0000000000000001: n9715_o = n9714_o;
      default: n9715_o = n9714_o;
    endcase
  assign n9716_o = sndopc[7];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9717_o = n9716_o;
      16'b0100000000000000: n9717_o = n9716_o;
      16'b0010000000000000: n9717_o = n9716_o;
      16'b0001000000000000: n9717_o = n9716_o;
      16'b0000100000000000: n9717_o = n9716_o;
      16'b0000010000000000: n9717_o = n9716_o;
      16'b0000001000000000: n9717_o = n9716_o;
      16'b0000000100000000: n9717_o = n9716_o;
      16'b0000000010000000: n9717_o = 1'b0;
      16'b0000000001000000: n9717_o = n9716_o;
      16'b0000000000100000: n9717_o = n9716_o;
      16'b0000000000010000: n9717_o = n9716_o;
      16'b0000000000001000: n9717_o = n9716_o;
      16'b0000000000000100: n9717_o = n9716_o;
      16'b0000000000000010: n9717_o = n9716_o;
      16'b0000000000000001: n9717_o = n9716_o;
      default: n9717_o = n9716_o;
    endcase
  assign n9718_o = sndopc[8];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9719_o = n9718_o;
      16'b0100000000000000: n9719_o = n9718_o;
      16'b0010000000000000: n9719_o = n9718_o;
      16'b0001000000000000: n9719_o = n9718_o;
      16'b0000100000000000: n9719_o = n9718_o;
      16'b0000010000000000: n9719_o = n9718_o;
      16'b0000001000000000: n9719_o = n9718_o;
      16'b0000000100000000: n9719_o = 1'b0;
      16'b0000000010000000: n9719_o = n9718_o;
      16'b0000000001000000: n9719_o = n9718_o;
      16'b0000000000100000: n9719_o = n9718_o;
      16'b0000000000010000: n9719_o = n9718_o;
      16'b0000000000001000: n9719_o = n9718_o;
      16'b0000000000000100: n9719_o = n9718_o;
      16'b0000000000000010: n9719_o = n9718_o;
      16'b0000000000000001: n9719_o = n9718_o;
      default: n9719_o = n9718_o;
    endcase
  assign n9720_o = sndopc[9];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9721_o = n9720_o;
      16'b0100000000000000: n9721_o = n9720_o;
      16'b0010000000000000: n9721_o = n9720_o;
      16'b0001000000000000: n9721_o = n9720_o;
      16'b0000100000000000: n9721_o = n9720_o;
      16'b0000010000000000: n9721_o = n9720_o;
      16'b0000001000000000: n9721_o = 1'b0;
      16'b0000000100000000: n9721_o = n9720_o;
      16'b0000000010000000: n9721_o = n9720_o;
      16'b0000000001000000: n9721_o = n9720_o;
      16'b0000000000100000: n9721_o = n9720_o;
      16'b0000000000010000: n9721_o = n9720_o;
      16'b0000000000001000: n9721_o = n9720_o;
      16'b0000000000000100: n9721_o = n9720_o;
      16'b0000000000000010: n9721_o = n9720_o;
      16'b0000000000000001: n9721_o = n9720_o;
      default: n9721_o = n9720_o;
    endcase
  assign n9722_o = sndopc[10];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9723_o = n9722_o;
      16'b0100000000000000: n9723_o = n9722_o;
      16'b0010000000000000: n9723_o = n9722_o;
      16'b0001000000000000: n9723_o = n9722_o;
      16'b0000100000000000: n9723_o = n9722_o;
      16'b0000010000000000: n9723_o = 1'b0;
      16'b0000001000000000: n9723_o = n9722_o;
      16'b0000000100000000: n9723_o = n9722_o;
      16'b0000000010000000: n9723_o = n9722_o;
      16'b0000000001000000: n9723_o = n9722_o;
      16'b0000000000100000: n9723_o = n9722_o;
      16'b0000000000010000: n9723_o = n9722_o;
      16'b0000000000001000: n9723_o = n9722_o;
      16'b0000000000000100: n9723_o = n9722_o;
      16'b0000000000000010: n9723_o = n9722_o;
      16'b0000000000000001: n9723_o = n9722_o;
      default: n9723_o = n9722_o;
    endcase
  assign n9724_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9725_o = n9724_o;
      16'b0100000000000000: n9725_o = n9724_o;
      16'b0010000000000000: n9725_o = n9724_o;
      16'b0001000000000000: n9725_o = n9724_o;
      16'b0000100000000000: n9725_o = 1'b0;
      16'b0000010000000000: n9725_o = n9724_o;
      16'b0000001000000000: n9725_o = n9724_o;
      16'b0000000100000000: n9725_o = n9724_o;
      16'b0000000010000000: n9725_o = n9724_o;
      16'b0000000001000000: n9725_o = n9724_o;
      16'b0000000000100000: n9725_o = n9724_o;
      16'b0000000000010000: n9725_o = n9724_o;
      16'b0000000000001000: n9725_o = n9724_o;
      16'b0000000000000100: n9725_o = n9724_o;
      16'b0000000000000010: n9725_o = n9724_o;
      16'b0000000000000001: n9725_o = n9724_o;
      default: n9725_o = n9724_o;
    endcase
  assign n9726_o = sndopc[12];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9727_o = n9726_o;
      16'b0100000000000000: n9727_o = n9726_o;
      16'b0010000000000000: n9727_o = n9726_o;
      16'b0001000000000000: n9727_o = 1'b0;
      16'b0000100000000000: n9727_o = n9726_o;
      16'b0000010000000000: n9727_o = n9726_o;
      16'b0000001000000000: n9727_o = n9726_o;
      16'b0000000100000000: n9727_o = n9726_o;
      16'b0000000010000000: n9727_o = n9726_o;
      16'b0000000001000000: n9727_o = n9726_o;
      16'b0000000000100000: n9727_o = n9726_o;
      16'b0000000000010000: n9727_o = n9726_o;
      16'b0000000000001000: n9727_o = n9726_o;
      16'b0000000000000100: n9727_o = n9726_o;
      16'b0000000000000010: n9727_o = n9726_o;
      16'b0000000000000001: n9727_o = n9726_o;
      default: n9727_o = n9726_o;
    endcase
  assign n9728_o = sndopc[13];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9729_o = n9728_o;
      16'b0100000000000000: n9729_o = n9728_o;
      16'b0010000000000000: n9729_o = 1'b0;
      16'b0001000000000000: n9729_o = n9728_o;
      16'b0000100000000000: n9729_o = n9728_o;
      16'b0000010000000000: n9729_o = n9728_o;
      16'b0000001000000000: n9729_o = n9728_o;
      16'b0000000100000000: n9729_o = n9728_o;
      16'b0000000010000000: n9729_o = n9728_o;
      16'b0000000001000000: n9729_o = n9728_o;
      16'b0000000000100000: n9729_o = n9728_o;
      16'b0000000000010000: n9729_o = n9728_o;
      16'b0000000000001000: n9729_o = n9728_o;
      16'b0000000000000100: n9729_o = n9728_o;
      16'b0000000000000010: n9729_o = n9728_o;
      16'b0000000000000001: n9729_o = n9728_o;
      default: n9729_o = n9728_o;
    endcase
  assign n9730_o = sndopc[14];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9731_o = n9730_o;
      16'b0100000000000000: n9731_o = 1'b0;
      16'b0010000000000000: n9731_o = n9730_o;
      16'b0001000000000000: n9731_o = n9730_o;
      16'b0000100000000000: n9731_o = n9730_o;
      16'b0000010000000000: n9731_o = n9730_o;
      16'b0000001000000000: n9731_o = n9730_o;
      16'b0000000100000000: n9731_o = n9730_o;
      16'b0000000010000000: n9731_o = n9730_o;
      16'b0000000001000000: n9731_o = n9730_o;
      16'b0000000000100000: n9731_o = n9730_o;
      16'b0000000000010000: n9731_o = n9730_o;
      16'b0000000000001000: n9731_o = n9730_o;
      16'b0000000000000100: n9731_o = n9730_o;
      16'b0000000000000010: n9731_o = n9730_o;
      16'b0000000000000001: n9731_o = n9730_o;
      default: n9731_o = n9730_o;
    endcase
  assign n9732_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9701_o)
      16'b1000000000000000: n9733_o = 1'b0;
      16'b0100000000000000: n9733_o = n9732_o;
      16'b0010000000000000: n9733_o = n9732_o;
      16'b0001000000000000: n9733_o = n9732_o;
      16'b0000100000000000: n9733_o = n9732_o;
      16'b0000010000000000: n9733_o = n9732_o;
      16'b0000001000000000: n9733_o = n9732_o;
      16'b0000000100000000: n9733_o = n9732_o;
      16'b0000000010000000: n9733_o = n9732_o;
      16'b0000000001000000: n9733_o = n9732_o;
      16'b0000000000100000: n9733_o = n9732_o;
      16'b0000000000010000: n9733_o = n9732_o;
      16'b0000000000001000: n9733_o = n9732_o;
      16'b0000000000000100: n9733_o = n9732_o;
      16'b0000000000000010: n9733_o = n9732_o;
      16'b0000000000000001: n9733_o = n9732_o;
      default: n9733_o = n9732_o;
    endcase
  assign n9734_o = {n9733_o, n9731_o, n9729_o, n9727_o, n9725_o, n9723_o, n9721_o, n9719_o, n9717_o, n9715_o, n9713_o, n9711_o, n9709_o, n9707_o, n9705_o, n9703_o};
  /* TG68KdotC_Kernel.vhd:4115:33  */
  assign n9735_o = n9652_o ? n9734_o : sndopc;
  /* TG68KdotC_Kernel.vhd:4113:33  */
  assign n9736_o = decodeopc ? n9649_o : n9735_o;
  /* TG68KdotC_Kernel.vhd:4144:26  */
  assign n9744_o = sndopc[3:0];
  /* TG68KdotC_Kernel.vhd:4144:38  */
  assign n9746_o = n9744_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4145:34  */
  assign n9747_o = sndopc[7:4];
  /* TG68KdotC_Kernel.vhd:4145:46  */
  assign n9749_o = n9747_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4147:42  */
  assign n9751_o = sndopc[11:8];
  /* TG68KdotC_Kernel.vhd:4147:55  */
  assign n9753_o = n9751_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4148:50  */
  assign n9754_o = sndopc[15:12];
  /* TG68KdotC_Kernel.vhd:4148:64  */
  assign n9756_o = n9754_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4148:41  */
  assign n9759_o = n9756_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:4152:60  */
  assign n9761_o = sndopc[15:12];
  /* TG68KdotC_Kernel.vhd:4154:60  */
  assign n9762_o = sndopc[11:8];
  /* TG68KdotC_Kernel.vhd:4147:33  */
  assign n9764_o = n9753_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:4147:33  */
  assign n9765_o = n9753_o ? n9761_o : n9762_o;
  /* TG68KdotC_Kernel.vhd:4147:33  */
  assign n9767_o = n9753_o ? n9759_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4157:52  */
  assign n9768_o = sndopc[7:4];
  assign n9770_o = {1'b1, n9764_o};
  assign n9771_o = n9770_o[0];
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9772_o = n9749_o ? n9771_o : 1'b1;
  assign n9773_o = n9770_o[1];
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9775_o = n9749_o ? n9773_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9776_o = n9749_o ? n9765_o : n9768_o;
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9778_o = n9749_o ? n9767_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4161:44  */
  assign n9779_o = sndopc[3:0];
  assign n9780_o = {n9775_o, n9772_o};
  /* TG68KdotC_Kernel.vhd:4144:17  */
  assign n9782_o = n9746_o ? n9780_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:4144:17  */
  assign n9785_o = n9746_o ? n9776_o : n9779_o;
  /* TG68KdotC_Kernel.vhd:4144:17  */
  assign n9787_o = n9746_o ? n9778_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4163:29  */
  assign n9789_o = movem_mux[1:0];
  /* TG68KdotC_Kernel.vhd:4163:41  */
  assign n9791_o = n9789_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:4165:37  */
  assign n9793_o = movem_mux[2];
  /* TG68KdotC_Kernel.vhd:4165:40  */
  assign n9794_o = ~n9793_o;
  assign n9796_o = n9783_o[0];
  /* TG68KdotC_Kernel.vhd:4165:25  */
  assign n9797_o = n9794_o ? 1'b1 : n9796_o;
  /* TG68KdotC_Kernel.vhd:4169:37  */
  assign n9798_o = movem_mux[0];
  /* TG68KdotC_Kernel.vhd:4169:40  */
  assign n9799_o = ~n9798_o;
  assign n9801_o = n9783_o[0];
  /* TG68KdotC_Kernel.vhd:4169:25  */
  assign n9802_o = n9799_o ? 1'b1 : n9801_o;
  assign n9803_o = {1'b1, n9797_o};
  assign n9804_o = n9803_o[0];
  /* TG68KdotC_Kernel.vhd:4163:17  */
  assign n9805_o = n9791_o ? n9804_o : n9802_o;
  assign n9806_o = n9803_o[1];
  assign n9807_o = n9783_o[1];
  /* TG68KdotC_Kernel.vhd:4163:17  */
  assign n9808_o = n9791_o ? n9806_o : n9807_o;
  /* TG68KdotC_Kernel.vhd:464:17  */
  always @(posedge clk)
    n9811_q <= n125_o;
  /* TG68KdotC_Kernel.vhd:458:17  */
  assign n9812_o = clkena_in ? n106_o : syncreset;
  /* TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n102_o)
    if (n102_o)
      n9813_q <= 4'b0000;
    else
      n9813_q <= n9812_o;
  /* TG68KdotC_Kernel.vhd:458:17  */
  assign n9814_o = clkena_in ? n108_o : reset;
  /* TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n102_o)
    if (n102_o)
      n9815_q <= 1'b1;
    else
      n9815_q <= n9814_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9816_q <= n1512_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9817_o = n1062_o ? addr : tmp_tg68_pc;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9818_q <= n9817_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9819_o = n1063_o ? addr : memaddr;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9820_q <= n9819_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9821_q <= n1514_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9822_q <= n1515_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9823_q <= n1517_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9824_q <= n1519_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9825_q <= n1520_o;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  assign n9826_o = clkena_lw ? n9736_o : sndopc;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  always @(posedge clk)
    n9827_q <= n9826_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9828_q <= n1521_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9829_q <= n1522_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9830_q <= n1524_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9832_o = clkena_lw ? rf_source_addr : rf_source_addrd;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9833_q <= n9832_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9834_o = {n356_o, n335_o, n353_o};
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9837_o = clkena_lw ? rf_dest_addr : rdindex_a;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9838_q <= n9837_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9839_o = clkena_lw ? rf_source_addr : rdindex_b;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9840_q <= n9839_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9841_o = clkena_lw ? n291_o : wr_areg;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9842_q <= n9841_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9843_o = clkena_in ? n1049_o : memaddr_delta_rega;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9844_q <= n9843_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9845_o = clkena_in ? n1051_o : memaddr_delta_regb;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9846_q <= n9845_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9847_o = clkena_in ? n1054_o : use_base;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9848_q <= n9847_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9849_q <= n790_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  assign n9850_o = {n619_o, n626_o};
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9852_q <= n791_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9853_q <= n1525_o;
  assign n9855_o = {n987_o, n984_o};
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9856_q <= n1527_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9857_q <= n1528_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9858_q <= n793_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9859_q <= n1530_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9860_q <= n1532_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9861_q <= n795_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9862_q <= n1534_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9863_q <= n1536_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9864_q <= n1538_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9865_q <= n1884_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9866_q <= n796_o;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  assign n9867_o = clkena_lw ? n1647_o : exec_tas;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  always @(posedge clk)
    n9868_q <= n9867_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9869_q <= n1539_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9870_q <= n1541_o;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  assign n9871_o = clkena_lw ? n9648_o : movem_actiond;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  always @(posedge clk)
    n9872_q <= n9871_o;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  assign n9873_o = {n9782_o, n9808_o, n9805_o};
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9875_q <= n798_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9876_q <= n800_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9877_q <= n1543_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9878_q <= n1545_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9879_q <= n1547_o;
  /* TG68KdotC_Kernel.vhd:3254:17  */
  always @(posedge clk)
    n9880_q <= n8144_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9881_q <= n1548_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9882_q <= n1886_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9883_q <= n1550_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9884_q <= n801_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9885_q <= n1552_o;
  /* TG68KdotC_Kernel.vhd:876:17  */
  assign n9886_o = clkena_lw ? n913_o : trap_vector;
  /* TG68KdotC_Kernel.vhd:876:17  */
  always @(posedge clk)
    n9887_q <= n9886_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9888_o = n306_o ? reg_qa : usp;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9889_q <= n9888_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9890_q <= n1553_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9891_q <= n1554_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9892_q <= n1556_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9893_q <= n1888_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9894_q <= n1890_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9895_q <= n1558_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9896_q <= n803_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  assign n9897_o = {n169_o, n172_o};
  /* TG68KdotC_Kernel.vhd:484:17  */
  assign n9898_o = n176_o ? n181_o : bf_ext_in;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9899_q <= n9898_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9900_q <= n1560_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9901_q <= n1561_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9902_q <= n1562_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9903_q <= n1563_o;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  always @(posedge clk)
    n9904_q <= n1617_o;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9905_q <= n228_o;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9906_q <= n229_o;
  /* TG68KdotC_Kernel.vhd:484:17  */
  assign n9907_o = {n1744_o, n1741_o, n1747_o};
  assign n9908_o = {1'b0, n1691_o};
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9909_q <= n1564_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9910_q <= n1565_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  assign n9911_o = {1'b0, n1704_o};
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9912_q <= n1566_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9913_q <= n1567_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9914_q <= n9510_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9915_q <= n9512_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9916_q <= n9513_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9917_q <= n9514_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  assign n9918_o = {n9375_o, n9373_o, n9371_o, n9367_o, n9363_o, n9359_o, n9358_o, n7956_o, n7932_o, n9357_o, n9416_o, n9415_o, n9355_o, n9351_o, n7927_o, n9350_o, n9349_o, n9348_o, n9347_o, n9412_o, n9343_o, n9409_o, n9339_o, n9403_o, n9338_o, n9334_o, n9330_o, n9326_o, n9394_o, n9322_o, n9321_o, n9388_o, n9317_o, n9316_o, n9315_o, n7918_o, n2002_o, n9314_o, n9310_o, n9306_o, n9305_o, n9382_o, n9301_o, n9300_o, n7945_o, n7911_o, n9379_o, n9299_o, n9297_o, n9296_o, n9295_o, n7940_o, n9294_o, n9293_o, n9292_o, n9378_o, n7939_o, n9288_o};
  assign n9919_o = {n7981_o, n8000_o, n7979_o, n7999_o, n7977_o, n7997_o, n7975_o, n7995_o, n8133_o, n8043_o, n7993_o, n8132_o, n7991_o, n8131_o, n9426_o, n9425_o, n9427_o, n7967_o, n7987_o, n7965_o, n7985_o, n7963_o};
  /* TG68KdotC_Kernel.vhd:1260:17  */
  assign n9920_o = clkena_lw ? n1661_o : exec;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  always @(posedge clk)
    n9921_q <= n9920_o;
  /* TG68KdotC_Kernel.vhd:3254:17  */
  always @(posedge clk)
    n9922_q <= n8146_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9923_q <= n1882_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9924_q <= n1510_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  assign n9925_o = {n9923_q, n9924_q};
  /* TG68KdotC_Kernel.vhd:558:35  */
  reg [31:0] regfile[15:0] ; // memory
  initial begin
    regfile[15] = 32'b00000000000000000000000000000000;
    regfile[14] = 32'b00000000000000000000000000000000;
    regfile[13] = 32'b00000000000000000000000000000000;
    regfile[12] = 32'b00000000000000000000000000000000;
    regfile[11] = 32'b00000000000000000000000000000000;
    regfile[10] = 32'b00000000000000000000000000000000;
    regfile[9] = 32'b00000000000000000000000000000000;
    regfile[8] = 32'b00000000000000000000000000000000;
    regfile[7] = 32'b00000000000000000000000000000000;
    regfile[6] = 32'b00000000000000000000000000000000;
    regfile[5] = 32'b00000000000000000000000000000000;
    regfile[4] = 32'b00000000000000000000000000000000;
    regfile[3] = 32'b00000000000000000000000000000000;
    regfile[2] = 32'b00000000000000000000000000000000;
    regfile[1] = 32'b00000000000000000000000000000000;
    regfile[0] = 32'b00000000000000000000000000000000;
    end
  assign n9927_data = regfile[rdindex_b];
  assign n9928_data = regfile[rdindex_a];
  always @(posedge clk)
    if (n302_o)
      regfile[rdindex_a] <= regin;
  /* TG68KdotC_Kernel.vhd:559:35  */
  /* TG68KdotC_Kernel.vhd:558:35  */
  /* TG68KdotC_Kernel.vhd:567:49  */
endmodule

module tg68kdotc_verilog_wrapper
  (input  clk,
   input  nReset,
   input  clkena_in,
   input  [15:0] data_in,
   input  [2:0] IPL,
   input  IPL_autovector,
   input  berr,
   output [31:0] addr_out,
   output [2:0] FC,
   output [15:0] data_write,
   output [1:0] busstate,
   output nWr,
   output nUDS,
   output nLDS,
   output nResetOut,
   output skipFetch);
  wire [31:0] tg68kdotcinst_addr_out;
  wire [15:0] tg68kdotcinst_data_write;
  wire tg68kdotcinst_nwr;
  wire tg68kdotcinst_nuds;
  wire tg68kdotcinst_nlds;
  wire [1:0] tg68kdotcinst_busstate;
  wire tg68kdotcinst_longword;
  wire tg68kdotcinst_nresetout;
  wire [2:0] tg68kdotcinst_fc;
  wire tg68kdotcinst_clr_berr;
  wire tg68kdotcinst_skipfetch;
  wire [31:0] tg68kdotcinst_regin_out;
  wire [3:0] tg68kdotcinst_cacr_out;
  wire [31:0] tg68kdotcinst_vbr_out;
  localparam [1:0] n9_o = 2'b01;
  assign addr_out = tg68kdotcinst_addr_out;
  assign FC = tg68kdotcinst_fc;
  assign data_write = tg68kdotcinst_data_write;
  assign busstate = tg68kdotcinst_busstate;
  assign nWr = tg68kdotcinst_nwr;
  assign nUDS = tg68kdotcinst_nuds;
  assign nLDS = tg68kdotcinst_nlds;
  assign nResetOut = tg68kdotcinst_nresetout;
  assign skipFetch = tg68kdotcinst_skipfetch;
  /* tg68dotc_verilog_wrapper.vhd:28:3  */
  tg68kdotc_kernel_2_2_2_2_2_2_1_1 tg68kdotcinst (
    .clk(clk),
    .nreset(nReset),
    .clkena_in(clkena_in),
    .data_in(data_in),
    .ipl(IPL),
    .ipl_autovector(IPL_autovector),
    .berr(berr),
    .cpu(n9_o),
    .addr_out(tg68kdotcinst_addr_out),
    .data_write(tg68kdotcinst_data_write),
    .nwr(tg68kdotcinst_nwr),
    .nuds(tg68kdotcinst_nuds),
    .nlds(tg68kdotcinst_nlds),
    .busstate(tg68kdotcinst_busstate),
    .longword(),
    .nresetout(tg68kdotcinst_nresetout),
    .fc(tg68kdotcinst_fc),
    .clr_berr(),
    .skipfetch(tg68kdotcinst_skipfetch),
    .regin_out(),
    .cacr_out(),
    .vbr_out());
endmodule

